CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
30
9 Resistor~
219 249 284 0 3 5
0 2 13 -1
0
0 0 96 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
43129.6 1
0
7 Ground~
168 249 319 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3951 0 0
2
43129.6 0
0
2 +V
167 405 343 0 1 3
0 18
0
0 0 53360 0
3 12V
13 -3 34 5
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
5.89833e-315 0
0
4 LED~
171 471 412 0 2 2
10 4 6
0
0 0 112 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3780 0 0
2
43129.6 0
0
7 Ground~
168 471 507 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
43129.6 1
0
11 SPDT Relay~
176 361 399 0 12 18
0 18 18 4 9 8 0 0 0 0
1 0 1
0
0 0 4208 0
7 12VSPDT
14 15 63 23
4 RLY2
21 4 49 12
0
0
20 %D %1 %2 %3 %4 %5 %S
0
16 alias:XSPDTRELAY
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 512 1 0 0 0
3 RLY
9442 0 0
2
43129.6 2
0
2 +V
167 243 354 0 1 3
0 9
0
0 0 53360 0
3 12V
13 -10 34 -2
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9424 0 0
2
43129.6 3
0
7 Ground~
168 243 504 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9968 0 0
2
43129.6 4
0
12 NPN Trans:B~
219 238 464 0 3 7
0 8 7 2
0
0 0 80 0
6 2N2222
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 1 0 0
1 Q
9281 0 0
2
43129.6 5
0
6 Diode~
219 243 414 0 2 5
0 8 9
0
0 0 80 90
6 1N4007
12 0 54 8
2 D1
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8464 0 0
2
43129.6 6
0
8 SPDT PB~
217 122 127 0 10 18
0 11 11 3 0 0 0 0 0 0
1
0
0 0 4208 0
0
3 S11
-8 -15 13 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7168 0 0
2
43129.6 7
0
4 4017
219 228 183 0 14 29
0 2 2 13 17 16 15 14 11 19
20 21 22 23 24
0
0 0 4208 90
4 4017
-14 -60 14 -52
2 U1
62 0 76 8
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
3171 0 0
2
43129.6 8
0
14 NO PushButton~
191 150 70 0 2 5
0 2 14
0
0 0 4208 90
0
2 S1
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4139 0 0
2
43129.6 10
0
2 +V
167 524 16 0 1 3
0 12
0
0 0 53360 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
43129.6 11
0
14 NO PushButton~
191 202 70 0 2 5
0 2 15
0
0 0 4208 90
0
2 S2
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5283 0 0
2
43129.6 12
0
14 NO PushButton~
191 251 70 0 2 5
0 2 16
0
0 0 4208 90
0
2 S3
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6874 0 0
2
43129.6 13
0
14 NO PushButton~
191 308 68 0 2 5
0 2 17
0
0 0 4208 90
0
2 S4
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5305 0 0
2
43129.6 14
0
14 NO PushButton~
191 390 80 0 2 5
0 12 13
0
0 0 4208 90
0
2 S5
14 -5 28 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
34 0 0
2
43129.6 15
0
14 NO PushButton~
191 440 79 0 2 5
0 12 13
0
0 0 4208 90
0
2 S6
16 -4 30 4
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
969 0 0
2
43129.6 16
0
14 NO PushButton~
191 490 81 0 2 5
0 12 13
0
0 0 4208 90
0
2 S7
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8402 0 0
2
43129.6 17
0
14 NO PushButton~
191 546 80 0 2 5
0 12 13
0
0 0 4208 90
0
2 S8
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3751 0 0
2
43129.6 18
0
14 NO PushButton~
191 598 80 0 2 5
0 12 13
0
0 0 4208 90
0
2 S9
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4292 0 0
2
43129.6 19
0
14 NO PushButton~
191 654 80 0 2 5
0 12 13
0
0 0 4208 90
0
3 S10
12 -5 33 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6118 0 0
2
43129.6 20
0
7 Ground~
168 311 321 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
34 0 0
2
43129.6 21
0
7 Ground~
168 202 321 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
43129.6 22
0
4 LED~
171 20 192 0 2 2
10 11 2
0
0 0 112 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
319 0 0
2
43129.6 23
0
7 Ground~
168 20 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3976 0 0
2
43129.6 24
0
9 Resistor~
219 471 462 0 4 5
0 6 2 0 -1
0
0 0 112 270
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7634 0 0
2
43129.6 25
0
9 Resistor~
219 137 464 0 2 5
0 7 3
0
0 0 112 180
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
523 0 0
2
43129.6 26
0
9 Resistor~
219 311 286 0 3 5
0 2 13 -1
0
0 0 112 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6748 0 0
2
43129.6 27
0
39
2 2 0 0 0 0 0 12 1 0 0 2
249 221
249 266
1 1 2 0 0 16 0 1 2 0 0 2
249 302
249 313
3 2 3 0 0 4224 0 11 29 0 0 3
105 141
105 464
119 464
3 1 4 0 0 4224 0 6 4 0 0 3
375 388
471 388
471 402
1 2 18 0 0 8320 5 3 6 0 0 5
405 352
405 370
383 370
383 374
375 374
1 2 2 0 0 4096 0 5 28 0 0 2
471 501
471 480
1 2 6 0 0 4224 0 28 4 0 0 2
471 444
471 422
1 2 7 0 0 4224 0 29 9 0 0 2
155 464
220 464
0 5 8 0 0 4224 0 0 6 13 0 4
243 434
346 434
346 418
345 418
0 4 9 0 0 4224 0 0 6 11 0 3
243 367
345 367
345 394
1 2 9 0 0 0 0 7 10 0 0 2
243 363
243 404
1 3 2 0 0 0 0 8 9 0 0 2
243 498
243 482
1 1 8 0 0 0 0 10 9 0 0 2
243 424
243 446
2 1 11 0 0 4224 10 11 26 0 0 3
105 127
20 127
20 182
1 8 11 0 0 4224 0 11 12 0 0 3
144 127
240 127
240 157
1 2 2 0 0 4096 0 27 26 0 0 2
20 242
20 202
1 0 12 0 0 4096 0 14 0 0 30 2
524 25
524 44
1 1 2 0 0 4096 0 25 12 0 0 4
202 315
202 228
240 228
240 227
0 0 13 0 0 8320 0 0 0 22 23 3
311 249
398 249
398 107
0 0 2 0 0 8320 0 0 0 0 33 4
249 238
346 238
346 36
313 36
1 1 2 0 0 0 0 30 24 0 0 2
311 304
311 315
2 3 13 0 0 0 0 30 12 0 0 4
311 268
311 248
267 248
267 221
0 2 13 0 0 0 0 0 18 24 0 3
448 107
398 107
398 97
0 2 13 0 0 0 0 0 19 25 0 3
500 107
448 107
448 96
0 2 13 0 0 0 0 0 20 26 0 3
554 107
498 107
498 98
0 2 13 0 0 0 0 0 21 27 0 3
608 107
554 107
554 97
2 2 13 0 0 0 0 23 22 0 0 4
662 97
662 107
606 107
606 97
0 1 12 0 0 4096 0 0 23 29 0 3
606 44
662 44
662 63
0 1 12 0 0 0 0 0 22 30 0 3
550 44
606 44
606 63
0 1 12 0 0 4224 0 0 21 31 0 3
497 44
554 44
554 63
0 1 12 0 0 0 0 0 20 32 0 3
448 44
498 44
498 64
1 1 12 0 0 0 0 18 19 0 0 4
398 63
398 44
448 44
448 62
0 1 2 0 0 0 0 0 17 34 0 3
259 36
316 36
316 51
0 1 2 0 0 0 0 0 16 35 0 3
210 36
259 36
259 53
1 1 2 0 0 0 0 13 15 0 0 4
158 53
158 36
210 36
210 53
7 2 14 0 0 8320 0 12 13 0 0 4
249 157
249 105
158 105
158 87
6 2 15 0 0 4224 0 12 15 0 0 4
258 157
258 98
210 98
210 87
5 2 16 0 0 4224 0 12 16 0 0 4
267 157
267 95
259 95
259 87
4 2 17 0 0 4224 0 12 17 0 0 4
276 157
276 93
316 93
316 85
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
