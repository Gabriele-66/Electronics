CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
820 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
79
13 Logic Switch~
5 1230 225 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
3 V18
8 -10 29 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
5.89821e-315 5.45523e-315
0
13 Logic Switch~
5 745 218 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
2 V1
11 -10 25 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.89821e-315 0
0
13 Logic Switch~
5 265 204 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
43036.5 0
0
2 +V
167 1324 449 0 1 3
0 7
0
0 0 53360 90
3 10V
6 -2 27 6
3 V17
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
961 0 0
2
5.89821e-315 5.45264e-315
0
7 Ground~
168 1457 446 0 1 3
0 2
0
0 0 53360 90
0
5 GND27
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
5.89821e-315 5.45005e-315
0
12 SPST Switch~
165 1405 447 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
6 reset2
-37 5 5 13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3409 0 0
2
5.89821e-315 5.44746e-315
0
5 4071~
219 1379 377 0 3 22
0 8 2 9
0
0 0 112 90
4 4071
-7 -24 21 -16
4 U10D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
3951 0 0
2
5.89821e-315 5.44487e-315
0
5 4081~
219 1282 260 0 3 22
0 12 13 11
0
0 0 112 270
4 4081
-7 -24 21 -16
4 U16B
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
8885 0 0
2
5.89821e-315 5.44228e-315
0
5 4081~
219 1020 266 0 3 22
0 14 15 10
0
0 0 112 270
4 4081
-7 -24 21 -16
4 U16A
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3780 0 0
2
5.89821e-315 5.43969e-315
0
5 4081~
219 1306 410 0 3 22
0 11 10 8
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U5D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
9265 0 0
2
5.89821e-315 5.4371e-315
0
7 Ground~
168 1411 311 0 1 3
0 2
0
0 0 53360 0
0
5 GND26
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9442 0 0
2
5.89821e-315 5.43192e-315
0
7 Ground~
168 1350 308 0 1 3
0 2
0
0 0 53360 0
0
5 GND25
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9424 0 0
2
5.89821e-315 5.42933e-315
0
7 Ground~
168 1138 310 0 1 3
0 2
0
0 0 53360 0
0
5 GND24
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9968 0 0
2
5.89821e-315 5.42414e-315
0
7 Ground~
168 1061 328 0 1 3
0 2
0
0 0 53360 0
0
5 GND23
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
5.89821e-315 5.41896e-315
0
2 +V
167 1074 320 0 1 3
0 17
0
0 0 53360 180
3 10V
6 -2 27 6
3 V15
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
5.89821e-315 5.41378e-315
0
9 CC 7-Seg~
183 1088 72 0 17 19
10 38 37 36 32 35 34 33 105 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7168 0 0
2
5.89821e-315 5.4086e-315
0
7 Ground~
168 1097 224 0 1 3
0 2
0
0 0 53360 0
0
5 GND22
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.89821e-315 5.40342e-315
0
2 +V
167 1383 223 0 1 3
0 19
0
0 0 53360 180
3 10V
6 -2 27 6
3 V14
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89821e-315 5.39824e-315
0
2 +V
167 1106 223 0 1 3
0 20
0
0 0 53360 180
3 10V
6 -2 27 6
3 V13
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89821e-315 5.39306e-315
0
7 Ground~
168 1374 226 0 1 3
0 2
0
0 0 53360 0
0
5 GND21
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5283 0 0
2
5.89821e-315 5.38788e-315
0
9 CC 7-Seg~
183 1365 74 0 17 19
10 29 28 27 23 26 25 24 106 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6874 0 0
2
5.89821e-315 5.37752e-315
0
4 4511
219 1365 178 0 20 29
0 13 22 21 12 2 19 18 24 25
26 23 27 28 29 0 0 0 0 0
9
0
0 0 4336 90
4 4511
-14 -60 14 -52
3 U15
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
5305 0 0
2
5.89821e-315 5.36716e-315
0
4 4029
219 1376 266 0 20 29
0 2 2 2 2 9 3 2 2 2
16 12 21 22 13 0 0 0 0 0
9
0
0 0 4336 90
4 4029
-14 -60 14 -52
3 U14
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
5.89821e-315 5.3568e-315
0
7 Ground~
168 1323 57 0 1 3
0 2
0
0 0 53360 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
969 0 0
2
5.89821e-315 5.34643e-315
0
7 Ground~
168 1129 49 0 1 3
0 2
0
0 0 53360 0
0
5 GND19
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8402 0 0
2
5.89821e-315 5.32571e-315
0
4 4029
219 1099 267 0 20 29
0 2 17 17 2 9 3 16 2 2
5 14 30 31 15 0 0 0 0 0
2
0
0 0 4336 90
4 4029
-14 -60 14 -52
3 U13
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
3751 0 0
2
5.89821e-315 5.30499e-315
0
4 4511
219 1088 179 0 20 29
0 15 31 30 14 2 20 18 33 34
35 32 36 37 38 0 0 0 0 0
2
0
0 0 4336 90
4 4511
-14 -60 14 -52
3 U12
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4292 0 0
2
5.89821e-315 5.26354e-315
0
4 4511
219 603 172 0 20 29
0 48 64 63 47 2 53 51 66 67
68 65 69 70 71 0 0 0 0 0
5
0
0 0 4336 90
4 4511
-14 -60 14 -52
3 U11
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6118 0 0
2
5.89821e-315 5.45264e-315
0
4 4029
219 614 260 0 20 29
0 2 50 50 2 42 3 49 2 2
4 47 63 64 48 0 0 0 0 0
5
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U9
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
5.89821e-315 5.45005e-315
0
7 Ground~
168 644 42 0 1 3
0 2
0
0 0 53360 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
5.89821e-315 5.44746e-315
0
7 Ground~
168 838 50 0 1 3
0 2
0
0 0 53360 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
319 0 0
2
5.89821e-315 5.44487e-315
0
4 4029
219 891 259 0 20 29
0 2 2 2 2 42 3 5 2 2
49 45 54 55 46 0 0 0 0 0
7
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
3976 0 0
2
5.89821e-315 5.44228e-315
0
4 4511
219 880 171 0 20 29
0 46 55 54 45 2 52 51 57 58
59 56 60 61 62 0 0 0 0 0
7
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U7
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7634 0 0
2
5.89821e-315 5.43969e-315
0
9 CC 7-Seg~
183 880 67 0 17 19
10 62 61 60 56 59 58 57 107 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
523 0 0
2
5.89821e-315 5.4371e-315
0
7 Ground~
168 889 219 0 1 3
0 2
0
0 0 53360 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6748 0 0
2
5.89821e-315 5.43451e-315
0
2 +V
167 621 216 0 1 3
0 53
0
0 0 53360 180
3 10V
6 -2 27 6
3 V12
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6901 0 0
2
5.89821e-315 5.43192e-315
0
2 +V
167 898 216 0 1 3
0 52
0
0 0 53360 180
3 10V
6 -2 27 6
3 V11
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
842 0 0
2
5.89821e-315 5.42933e-315
0
7 Ground~
168 612 217 0 1 3
0 2
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3277 0 0
2
5.89821e-315 5.42414e-315
0
9 CC 7-Seg~
183 603 65 0 17 19
10 71 70 69 65 68 67 66 108 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4212 0 0
2
5.89821e-315 5.41896e-315
0
2 +V
167 589 313 0 1 3
0 50
0
0 0 53360 180
3 10V
6 -2 27 6
2 V9
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4720 0 0
2
5.89821e-315 5.41378e-315
0
7 Ground~
168 576 321 0 1 3
0 2
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5551 0 0
2
5.89821e-315 5.4086e-315
0
7 Ground~
168 654 301 0 1 3
0 2
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
5.89821e-315 5.40342e-315
0
7 Ground~
168 865 301 0 1 3
0 2
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8745 0 0
2
5.89821e-315 5.39824e-315
0
7 Ground~
168 934 306 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9592 0 0
2
5.89821e-315 5.39306e-315
0
7 Pulser~
4 730 504 0 10 12
0 109 110 3 111 0 0 5 5 6
7
0
0 0 5168 0
0
2 V4
-8 -28 6 -20
15 automatic clock
-52 -28 53 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8748 0 0
2
5.89821e-315 5.38788e-315
0
5 4081~
219 821 403 0 3 22
0 44 43 41
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7168 0 0
2
5.89821e-315 5.37752e-315
0
5 4081~
219 535 259 0 3 22
0 47 48 43
0
0 0 112 270
4 4081
-7 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
631 0 0
2
5.89821e-315 5.36716e-315
0
5 4081~
219 797 253 0 3 22
0 45 46 44
0
0 0 112 270
4 4081
-7 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9466 0 0
2
5.89821e-315 5.3568e-315
0
5 4071~
219 894 370 0 3 22
0 41 2 42
0
0 0 112 90
4 4071
-7 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
3266 0 0
2
5.89821e-315 5.34643e-315
0
12 SPST Switch~
165 920 440 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
6 reset1
-37 5 5 13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7693 0 0
2
5.89821e-315 5.32571e-315
0
7 Ground~
168 972 439 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3723 0 0
2
5.89821e-315 5.30499e-315
0
2 +V
167 839 442 0 1 3
0 40
0
0 0 53360 90
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3440 0 0
2
5.89821e-315 5.26354e-315
0
2 +V
167 359 428 0 1 3
0 73
0
0 0 53360 90
3 10V
6 -2 27 6
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6263 0 0
2
43036.5 1
0
7 Ground~
168 492 425 0 1 3
0 2
0
0 0 53360 90
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4900 0 0
2
43036.5 2
0
12 SPST Switch~
165 440 426 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
5 reset
-34 5 1 13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8783 0 0
2
43036.5 3
0
5 4071~
219 414 356 0 3 22
0 74 2 75
0
0 0 112 90
4 4071
-7 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
3221 0 0
2
43036.5 4
0
5 4081~
219 317 239 0 3 22
0 78 79 77
0
0 0 112 270
4 4081
-7 -24 21 -16
3 U6D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3215 0 0
2
43036.5 5
0
5 4081~
219 55 245 0 3 22
0 80 81 76
0
0 0 112 270
4 4081
-7 -24 21 -16
3 U6C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7903 0 0
2
43036.5 6
0
5 4081~
219 341 389 0 3 22
0 77 76 74
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
7121 0 0
2
43036.5 7
0
7 Ground~
168 454 292 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4484 0 0
2
5.89821e-315 0
0
7 Ground~
168 385 287 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5996 0 0
2
5.89821e-315 5.26354e-315
0
7 Ground~
168 173 289 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7804 0 0
2
5.89821e-315 5.30499e-315
0
7 Ground~
168 96 307 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5523 0 0
2
5.89821e-315 5.32571e-315
0
2 +V
167 109 299 0 1 3
0 83
0
0 0 53360 180
3 10V
6 -2 27 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3330 0 0
2
5.89821e-315 5.34643e-315
0
9 CC 7-Seg~
183 123 51 0 17 19
10 104 103 102 98 101 100 99 112 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3465 0 0
2
43036.5 8
0
7 Ground~
168 132 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8396 0 0
2
43036.5 9
0
2 +V
167 418 202 0 1 3
0 85
0
0 0 53360 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3685 0 0
2
43036.5 10
0
2 +V
167 141 202 0 1 3
0 86
0
0 0 53360 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7849 0 0
2
43036.5 11
0
7 Ground~
168 409 205 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6343 0 0
2
43036.5 12
0
9 CC 7-Seg~
183 400 53 0 17 19
10 95 94 93 89 92 91 90 113 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7376 0 0
2
43036.5 13
0
4 4511
219 400 157 0 14 29
0 79 88 87 78 2 85 84 90 91
92 89 93 94 95
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
9156 0 0
2
43036.5 14
0
4 4029
219 411 245 0 14 29
0 2 2 2 2 75 3 4 2 2
82 78 87 88 79
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
5776 0 0
2
43036.5 15
0
7 Ground~
168 358 36 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7207 0 0
2
43036.5 16
0
7 Ground~
168 164 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4459 0 0
2
43036.5 17
0
4 4029
219 134 246 0 20 29
0 2 83 83 2 75 3 82 2 2
114 80 96 97 81 0 0 0 0 0
6
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 512 1 0 0 0
1 U
3760 0 0
2
5.89821e-315 5.3568e-315
0
4 4511
219 123 158 0 20 29
0 81 97 96 80 2 86 84 99 100
101 98 102 103 104 0 0 0 0 0
6
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
754 0 0
2
5.89821e-315 5.36716e-315
0
13 SemiResistor~
219 1362 447 0 4 5
0 2 7 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R2
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9767 0 0
2
5.89821e-315 0
0
13 SemiResistor~
219 877 440 0 4 5
0 2 40 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R1
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7978 0 0
2
5.89821e-315 5.45523e-315
0
13 SemiResistor~
219 397 426 0 4 5
0 2 73 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R6
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3142 0 0
2
43036.5 18
0
177
0 0 3 0 0 4096 0 0 0 2 24 3
769 457
1248 457
1248 335
0 0 3 0 0 8320 0 0 0 138 76 3
272 314
272 457
769 457
10 7 4 0 0 4224 0 29 72 0 0 5
621 224
486 224
486 312
436 312
436 285
10 7 5 0 0 4224 0 26 32 0 0 5
1106 231
973 231
973 302
916 302
916 299
8 9 2 0 0 4096 0 32 32 0 0 2
925 293
934 293
2 2 2 0 0 4224 6 7 6 0 0 3
1391 393
1391 447
1388 447
1 1 2 0 0 4096 0 5 6 0 0 2
1450 447
1422 447
2 1 2 0 0 0 6 6 77 0 0 2
1388 447
1380 447
2 1 7 0 0 4224 0 77 4 0 0 2
1344 447
1335 447
3 1 8 0 0 4224 0 10 7 0 0 3
1327 410
1373 410
1373 393
3 0 9 0 0 4096 0 7 0 0 18 2
1382 347
1382 348
3 2 10 0 0 8320 0 9 10 0 0 3
1018 289
1018 419
1282 419
3 1 11 0 0 4224 0 8 10 0 0 3
1280 283
1280 401
1282 401
1 0 12 0 0 8320 0 8 0 0 41 3
1289 238
1289 219
1365 219
2 0 13 0 0 8320 0 8 0 0 44 3
1271 238
1271 214
1338 214
1 0 14 0 0 8320 0 9 0 0 53 3
1027 244
1027 221
1088 221
2 0 15 0 0 8320 0 9 0 0 56 3
1009 244
1009 206
1061 206
5 5 9 0 0 8320 0 26 23 0 0 4
1106 301
1106 348
1383 348
1383 300
9 1 2 0 0 0 0 26 13 0 0 3
1142 301
1142 304
1138 304
8 1 2 0 0 0 0 26 13 0 0 3
1133 301
1133 304
1138 304
9 1 2 0 0 0 0 23 11 0 0 3
1419 300
1419 305
1411 305
8 1 2 0 0 0 0 23 11 0 0 3
1410 300
1410 305
1411 305
7 1 2 0 0 0 0 23 11 0 0 3
1401 306
1401 305
1411 305
6 6 3 0 0 0 0 26 23 0 0 4
1115 301
1115 335
1392 335
1392 300
7 10 16 0 0 8320 0 26 23 0 0 5
1124 307
1124 324
1436 324
1436 230
1383 230
1 4 2 0 0 0 0 14 26 0 0 3
1061 322
1088 322
1088 301
1 1 2 0 0 0 0 26 14 0 0 2
1061 301
1061 322
1 0 17 0 0 4096 0 15 0 0 29 2
1074 305
1074 301
2 3 17 0 0 4224 0 26 26 0 0 2
1070 301
1079 301
1 0 2 0 0 0 0 12 0 0 32 3
1350 302
1350 300
1351 300
4 3 2 0 0 0 0 23 23 0 0 2
1365 300
1356 300
3 2 2 0 0 0 0 23 23 0 0 2
1356 300
1347 300
1 2 2 0 0 0 0 23 23 0 0 2
1338 300
1347 300
1 0 18 0 0 12288 0 1 0 0 35 6
1231 212
1231 213
1231 213
1231 201
1230 201
1230 202
7 7 18 0 0 4224 0 27 22 0 0 3
1115 202
1392 202
1392 201
6 1 19 0 0 4224 0 22 18 0 0 4
1383 201
1383 209
1383 209
1383 208
5 1 2 0 0 0 0 22 20 0 0 2
1374 201
1374 220
6 1 20 0 0 4224 0 27 19 0 0 4
1106 202
1106 210
1106 210
1106 208
5 1 2 0 0 0 0 27 17 0 0 2
1097 202
1097 218
9 1 2 0 0 8320 0 21 24 0 0 4
1365 32
1365 28
1323 28
1323 51
4 11 12 0 0 0 0 22 23 0 0 2
1365 195
1365 236
3 12 21 0 0 4224 0 22 23 0 0 2
1356 195
1356 236
2 13 22 0 0 4224 0 22 23 0 0 2
1347 195
1347 236
1 14 13 0 0 0 0 22 23 0 0 2
1338 195
1338 236
4 11 23 0 0 4224 0 21 22 0 0 3
1362 110
1362 131
1365 131
7 8 24 0 0 4224 0 21 22 0 0 4
1380 110
1380 124
1392 124
1392 131
6 9 25 0 0 4224 0 21 22 0 0 4
1374 110
1374 129
1383 129
1383 131
5 10 26 0 0 4224 0 21 22 0 0 3
1368 110
1368 131
1374 131
3 12 27 0 0 4224 0 21 22 0 0 2
1356 110
1356 131
2 13 28 0 0 4224 0 21 22 0 0 3
1350 110
1350 131
1347 131
1 14 29 0 0 4224 0 21 22 0 0 3
1344 110
1344 131
1338 131
9 1 2 0 0 0 0 16 25 0 0 4
1088 30
1088 27
1129 27
1129 43
4 11 14 0 0 0 0 27 26 0 0 2
1088 196
1088 237
3 12 30 0 0 4224 0 27 26 0 0 2
1079 196
1079 237
2 13 31 0 0 4224 0 27 26 0 0 2
1070 196
1070 237
1 14 15 0 0 0 0 27 26 0 0 2
1061 196
1061 237
4 11 32 0 0 4224 0 16 27 0 0 4
1085 108
1085 133
1088 133
1088 132
7 8 33 0 0 4224 0 16 27 0 0 4
1103 108
1103 123
1115 123
1115 132
6 9 34 0 0 4224 0 16 27 0 0 4
1097 108
1097 128
1106 128
1106 132
5 10 35 0 0 4224 0 16 27 0 0 4
1091 108
1091 133
1097 133
1097 132
3 12 36 0 0 4224 0 16 27 0 0 2
1079 108
1079 132
2 13 37 0 0 4224 0 16 27 0 0 4
1073 108
1073 133
1070 133
1070 132
1 14 38 0 0 4224 0 16 27 0 0 4
1067 108
1067 133
1061 133
1061 132
2 2 2 0 0 4224 39 49 50 0 0 3
906 386
906 440
903 440
1 1 2 0 0 0 0 51 50 0 0 2
965 440
937 440
2 1 2 0 0 0 39 50 78 0 0 2
903 440
895 440
2 1 40 0 0 4224 0 78 52 0 0 2
859 440
850 440
3 1 41 0 0 4224 0 46 49 0 0 3
842 403
888 403
888 386
3 0 42 0 0 4096 0 49 0 0 77 2
897 340
897 341
3 2 43 0 0 8320 0 47 46 0 0 3
533 282
533 412
797 412
3 1 44 0 0 4224 0 48 46 0 0 3
795 276
795 394
797 394
1 0 45 0 0 8320 0 48 0 0 98 3
804 231
804 212
880 212
2 0 46 0 0 8320 0 48 0 0 101 3
786 231
786 207
853 207
1 0 47 0 0 8320 0 47 0 0 110 3
542 237
542 214
603 214
2 0 48 0 0 8320 0 47 0 0 113 3
524 237
524 199
576 199
3 0 3 0 0 0 0 45 0 0 81 3
754 495
769 495
769 328
5 5 42 0 0 8320 0 29 32 0 0 4
621 294
621 341
898 341
898 293
9 1 2 0 0 0 0 29 42 0 0 4
657 294
657 296
654 296
654 295
8 1 2 0 0 0 0 29 42 0 0 3
648 294
648 295
654 295
9 1 2 0 0 0 0 32 44 0 0 2
934 293
934 300
6 6 3 0 0 0 0 29 32 0 0 4
630 294
630 328
907 328
907 293
7 10 49 0 0 8320 0 29 32 0 0 5
639 300
639 317
951 317
951 223
898 223
1 4 2 0 0 0 0 41 29 0 0 3
576 315
603 315
603 294
1 1 2 0 0 0 0 29 41 0 0 2
576 294
576 315
1 0 50 0 0 4096 0 40 0 0 86 2
589 298
589 294
2 3 50 0 0 4224 0 29 29 0 0 2
585 294
594 294
1 0 2 0 0 0 0 43 0 0 89 3
865 295
865 293
866 293
4 3 2 0 0 0 0 32 32 0 0 2
880 293
871 293
3 2 2 0 0 0 0 32 32 0 0 2
871 293
862 293
1 2 2 0 0 0 0 32 32 0 0 2
853 293
862 293
1 0 51 0 0 12288 0 2 0 0 92 6
746 205
746 206
746 206
746 194
745 194
745 195
7 7 51 0 0 4224 0 28 33 0 0 3
630 195
907 195
907 194
6 1 52 0 0 4224 0 33 37 0 0 4
898 194
898 202
898 202
898 201
5 1 2 0 0 0 0 33 35 0 0 2
889 194
889 213
6 1 53 0 0 4224 0 28 36 0 0 4
621 195
621 203
621 203
621 201
5 1 2 0 0 0 0 28 38 0 0 2
612 195
612 211
9 1 2 0 0 0 0 34 31 0 0 4
880 25
880 21
838 21
838 44
4 11 45 0 0 0 0 33 32 0 0 2
880 188
880 229
3 12 54 0 0 4224 0 33 32 0 0 2
871 188
871 229
2 13 55 0 0 4224 0 33 32 0 0 2
862 188
862 229
1 14 46 0 0 0 0 33 32 0 0 2
853 188
853 229
4 11 56 0 0 4224 0 34 33 0 0 3
877 103
877 124
880 124
7 8 57 0 0 4224 0 34 33 0 0 4
895 103
895 117
907 117
907 124
6 9 58 0 0 4224 0 34 33 0 0 4
889 103
889 122
898 122
898 124
5 10 59 0 0 4224 0 34 33 0 0 3
883 103
883 124
889 124
3 12 60 0 0 4224 0 34 33 0 0 2
871 103
871 124
2 13 61 0 0 4224 0 34 33 0 0 3
865 103
865 124
862 124
1 14 62 0 0 4224 0 34 33 0 0 3
859 103
859 124
853 124
9 1 2 0 0 0 0 39 30 0 0 4
603 23
603 20
644 20
644 36
4 11 47 0 0 0 0 28 29 0 0 2
603 189
603 230
3 12 63 0 0 4224 0 28 29 0 0 2
594 189
594 230
2 13 64 0 0 4224 0 28 29 0 0 2
585 189
585 230
1 14 48 0 0 0 0 28 29 0 0 2
576 189
576 230
4 11 65 0 0 4224 0 39 28 0 0 4
600 101
600 126
603 126
603 125
7 8 66 0 0 4224 0 39 28 0 0 4
618 101
618 116
630 116
630 125
6 9 67 0 0 4224 0 39 28 0 0 4
612 101
612 121
621 121
621 125
5 10 68 0 0 4224 0 39 28 0 0 4
606 101
606 126
612 126
612 125
3 12 69 0 0 4224 0 39 28 0 0 2
594 101
594 125
2 13 70 0 0 4224 0 39 28 0 0 4
588 101
588 126
585 126
585 125
1 14 71 0 0 4224 0 39 28 0 0 4
582 101
582 126
576 126
576 125
2 2 2 0 0 4224 72 56 55 0 0 3
426 372
426 426
423 426
1 1 2 0 0 0 0 54 55 0 0 2
485 426
457 426
2 1 2 0 0 0 72 55 79 0 0 2
423 426
415 426
2 1 73 0 0 4224 0 79 53 0 0 2
379 426
370 426
3 1 74 0 0 4224 0 59 56 0 0 3
362 389
408 389
408 372
3 0 75 0 0 4096 0 56 0 0 133 2
417 326
417 327
3 2 76 0 0 8320 0 58 59 0 0 3
53 268
53 398
317 398
3 1 77 0 0 4224 0 57 59 0 0 3
315 262
315 380
317 380
1 0 78 0 0 8320 0 57 0 0 155 3
324 217
324 198
400 198
2 0 79 0 0 8320 0 57 0 0 158 3
306 217
306 193
373 193
1 0 80 0 0 8320 0 58 0 0 167 3
62 223
62 200
123 200
2 0 81 0 0 8320 0 58 0 0 170 3
44 223
44 185
96 185
5 5 75 0 0 8320 0 75 72 0 0 4
141 280
141 327
418 327
418 279
9 1 2 0 0 0 0 75 62 0 0 3
177 280
177 283
173 283
8 1 2 0 0 0 0 75 62 0 0 3
168 280
168 283
173 283
9 1 2 0 0 0 0 72 60 0 0 2
454 279
454 286
8 1 2 0 0 0 0 72 60 0 0 3
445 279
445 286
454 286
6 6 3 0 0 0 0 75 72 0 0 4
150 280
150 314
427 314
427 279
7 10 82 0 0 8320 0 75 72 0 0 5
159 286
159 303
471 303
471 209
418 209
1 4 2 0 0 0 0 63 75 0 0 3
96 301
123 301
123 280
1 1 2 0 0 0 0 75 63 0 0 2
96 280
96 301
1 0 83 0 0 4096 0 64 0 0 143 2
109 284
109 280
2 3 83 0 0 4224 0 75 75 0 0 2
105 280
114 280
1 0 2 0 0 0 0 61 0 0 146 3
385 281
385 279
386 279
4 3 2 0 0 0 0 72 72 0 0 2
400 279
391 279
3 2 2 0 0 0 0 72 72 0 0 2
391 279
382 279
1 2 2 0 0 0 0 72 72 0 0 2
373 279
382 279
1 0 84 0 0 12288 0 3 0 0 149 6
266 191
266 192
266 192
266 180
265 180
265 181
7 7 84 0 0 4224 0 76 71 0 0 3
150 181
427 181
427 180
6 1 85 0 0 4224 0 71 67 0 0 4
418 180
418 188
418 188
418 187
5 1 2 0 0 0 0 71 69 0 0 2
409 180
409 199
6 1 86 0 0 4224 0 76 68 0 0 4
141 181
141 189
141 189
141 187
5 1 2 0 0 0 0 76 66 0 0 2
132 181
132 197
9 1 2 0 0 0 0 70 73 0 0 4
400 11
400 7
358 7
358 30
4 11 78 0 0 0 0 71 72 0 0 2
400 174
400 215
3 12 87 0 0 4224 0 71 72 0 0 2
391 174
391 215
2 13 88 0 0 4224 0 71 72 0 0 2
382 174
382 215
1 14 79 0 0 0 0 71 72 0 0 2
373 174
373 215
4 11 89 0 0 4224 0 70 71 0 0 3
397 89
397 110
400 110
7 8 90 0 0 4224 0 70 71 0 0 4
415 89
415 103
427 103
427 110
6 9 91 0 0 4224 0 70 71 0 0 4
409 89
409 108
418 108
418 110
5 10 92 0 0 4224 0 70 71 0 0 3
403 89
403 110
409 110
3 12 93 0 0 4224 0 70 71 0 0 2
391 89
391 110
2 13 94 0 0 4224 0 70 71 0 0 3
385 89
385 110
382 110
1 14 95 0 0 4224 0 70 71 0 0 3
379 89
379 110
373 110
9 1 2 0 0 0 0 65 74 0 0 4
123 9
123 6
164 6
164 22
4 11 80 0 0 0 0 76 75 0 0 2
123 175
123 216
3 12 96 0 0 4224 0 76 75 0 0 2
114 175
114 216
2 13 97 0 0 4224 0 76 75 0 0 2
105 175
105 216
1 14 81 0 0 0 0 76 75 0 0 2
96 175
96 216
4 11 98 0 0 4224 0 65 76 0 0 4
120 87
120 112
123 112
123 111
7 8 99 0 0 4224 0 65 76 0 0 4
138 87
138 102
150 102
150 111
6 9 100 0 0 4224 0 65 76 0 0 4
132 87
132 107
141 107
141 111
5 10 101 0 0 4224 0 65 76 0 0 4
126 87
126 112
132 112
132 111
3 12 102 0 0 4224 0 65 76 0 0 2
114 87
114 111
2 13 103 0 0 4224 0 65 76 0 0 4
108 87
108 112
105 112
105 111
1 14 104 0 0 4224 0 65 76 0 0 4
102 87
102 112
96 112
96 111
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
