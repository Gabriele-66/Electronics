CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
46
12 PNP Trans:B~
219 609 71 0 3 7
0 6 14 13
0
0 0 832 692
5 BC327
-58 -15 -23 -7
2 Q2
-49 -27 -35 -19
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
113 0 0 0 1 0 0 0
1 Q
5130 0 0
2
43528.4 2
0
2 +V
167 614 33 0 1 3
0 13
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
43528.4 1
0
9 Resistor~
219 645 91 0 2 5
0 6 40
0
0 0 864 0
7 560 ohm
-24 -14 25 -6
2 R9
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 1 0 0 0
1 R
3124 0 0
2
43528.4 0
0
2 +V
167 605 282 0 1 3
0 7
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 V12
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3421 0 0
2
43528.4 8
0
12 PNP Trans:B~
219 601 317 0 3 7
0 26 8 7
0
0 0 320 692
5 BC327
2 -5 37 3
2 Q4
27 -10 41 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
113 0 0 512 1 0 0 0
1 Q
8157 0 0
2
43528.4 7
0
9 Resistor~
219 661 335 0 2 5
0 6 40
0
0 0 864 0
7 220 ohm
-24 -14 25 -6
3 R16
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 1 0 0 0
1 R
5572 0 0
2
43528.4 6
0
2 +V
167 545 259 0 1 3
0 4
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
43528.4 5
0
7 Ground~
168 454 354 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
43528.4 4
0
2 +V
167 454 289 0 1 3
0 11
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
43528.4 3
0
12 Comparator5~
219 454 320 0 5 11
0 12 9 2 11 5
0
0 0 320 692
5 LM339
5 -15 40 -7
2 U3
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 0 0 0
1 U
972 0 0
2
43528.4 2
0
9 Resistor~
219 545 292 0 4 5
0 5 4 0 1
0
0 0 864 90
3 22k
8 4 29 12
3 R14
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3472 0 0
2
43528.4 1
0
9 Resistor~
219 566 320 0 2 5
0 5 39
0
0 0 864 0
3 22k
-10 9 11 17
3 R15
-11 19 10 27
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 1 0 0 0
1 R
9998 0 0
2
43528.4 0
0
7 Ground~
168 465 238 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
43528.4 0
0
9 Resistor~
219 73 250 0 3 5
0 2 24 -1
0
0 0 864 90
4 270k
-33 1 -5 9
2 R3
-20 -9 -6 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
43528.4 45
0
9 Resistor~
219 44 211 0 2 5
0 3 24
0
0 0 864 0
2 1k
-7 7 7 15
2 R1
-7 -14 7 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
43528.4 44
0
9 Resistor~
219 163 314 0 3 5
0 2 20 -1
0
0 0 864 0
3 15k
-11 -14 10 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
43528.4 43
0
9 Resistor~
219 73 172 0 4 5
0 24 25 0 1
0
0 0 864 90
4 680k
-39 3 -11 11
2 R2
-20 -10 -6 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5616 0 0
2
43528.4 42
0
9 Resistor~
219 263 315 0 4 5
0 12 21 0 1
0
0 0 864 0
3 56k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
43528.4 41
0
9 Resistor~
219 218 314 0 2 5
0 20 12
0
0 0 864 0
3 22k
-11 -14 10 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
43528.4 40
0
9 Resistor~
219 414 183 0 4 5
0 17 16 0 1
0
0 0 864 90
4 330k
1 0 29 8
3 R10
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
43528.4 39
0
9 Resistor~
219 356 133 0 2 5
0 15 14
0
0 0 864 0
4 4.7k
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
43528.4 38
0
9 Resistor~
219 313 115 0 4 5
0 15 18 0 1
0
0 0 864 90
3 22k
5 0 26 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
43528.4 37
0
9 Resistor~
219 568 212 0 2 5
0 9 8
0
0 0 864 0
3 12k
-10 -14 11 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
43528.4 36
0
9 Resistor~
219 517 188 0 4 5
0 9 10 0 1
0
0 0 864 90
3 22k
8 0 29 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
43528.4 35
0
12 Comparator5~
219 259 133 0 5 11
0 24 20 23 2 15
0
0 0 320 0
5 LM339
5 -18 40 -10
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 0 0 0
1 U
9172 0 0
2
43528.4 31
0
12 Comparator5~
219 254 245 0 5 11
0 12 24 22 2 17
0
0 0 320 0
5 LM339
12 -16 47 -8
2 U2
4 -35 18 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 0 0 0
1 U
7100 0 0
2
43528.4 30
0
12 Comparator5~
219 465 212 0 5 11
0 17 12 2 19 9
0
0 0 320 692
5 LM339
8 -21 43 -13
2 U4
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 0 0 0
1 U
3820 0 0
2
43528.4 28
0
2 +V
167 93 88 0 1 3
0 25
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 Vcc
-11 -15 10 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
43528.4 27
0
2 +V
167 517 155 0 1 3
0 10
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
961 0 0
2
43528.4 26
0
2 +V
167 414 151 0 1 3
0 16
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3178 0 0
2
43528.4 25
0
2 +V
167 313 56 0 1 3
0 18
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V5
-7 -28 7 -20
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
43528.4 23
0
2 +V
167 465 169 0 1 3
0 19
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
43528.4 22
0
2 +V
167 613 130 0 1 3
0 7
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
43528.4 20
0
2 +V
167 254 216 0 1 3
0 22
0
0 0 53472 0
3 10V
-11 -15 10 -7
2 V9
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3780 0 0
2
43528.4 19
0
2 +V
167 306 306 0 1 3
0 21
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9265 0 0
2
43528.4 18
0
2 +V
167 259 98 0 1 3
0 23
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
43528.4 17
0
6 Diode~
219 109 177 0 2 5
0 24 25
0
0 0 832 90
6 1N4148
12 0 54 8
2 D1
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9424 0 0
2
43528.4 16
0
6 Diode~
219 109 251 0 2 5
0 2 24
0
0 0 832 90
6 1N4148
12 0 54 8
2 D2
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9968 0 0
2
43528.4 15
0
6 Diode~
219 336 205 0 2 5
0 17 15
0
0 0 320 180
6 1N4148
-21 -18 21 -10
2 D3
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9281 0 0
2
43528.4 14
0
11 Terminal:A~
194 20 211 0 1 3
0 3
0
0 0 57568 0
3 Vin
-10 -13 11 -5
2 J1
-7 -23 7 -15
0
4 Vin;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
8464 0 0
2
43528.4 13
0
7 Ground~
168 259 158 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
43528.4 12
0
7 Ground~
168 140 326 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
43528.4 11
0
7 Ground~
168 30 299 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4139 0 0
2
43528.4 10
0
7 Ground~
168 254 268 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
43528.4 8
0
12 PNP Trans:B~
219 608 176 0 3 7
0 26 8 7
0
0 0 320 692
5 BC327
6 -3 41 5
2 Q3
27 -10 41 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
113 0 0 512 1 0 0 0
1 Q
5283 0 0
2
43528.4 6
0
9 Resistor~
219 673 194 0 2 5
0 6 40
0
0 0 864 0
2 1k
-7 -14 7 -6
3 R13
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 1 0 0 0
1 R
6874 0 0
2
43528.4 3
0
51
1 1 6 0 0 0 0 3 1 0 0 3
627 91
614 91
614 89
1 3 13 0 0 0 0 2 1 0 0 2
614 42
614 53
2 0 0 0 0 0 0 10 0 0 15 5
436 326
426 326
426 256
517 256
517 212
0 0 0 0 0 0 0 0 0 25 5 2
236 286
415 286
2 1 0 0 0 0 0 27 10 0 0 4
447 218
415 218
415 314
436 314
2 2 0 0 0 0 0 5 12 0 0 3
583 317
583 320
584 320
1 1 0 0 0 0 0 6 5 0 0 2
643 335
606 335
1 3 7 0 0 0 0 4 5 0 0 4
605 291
605 296
606 296
606 299
1 2 4 0 0 0 0 7 11 0 0 2
545 268
545 274
1 0 5 0 0 0 0 11 0 0 11 2
545 310
545 320
1 5 5 0 0 0 0 12 10 0 0 2
548 320
472 320
1 3 2 0 0 0 0 8 10 0 0 2
454 348
454 333
1 4 11 0 0 0 0 9 10 0 0 2
454 298
454 307
1 3 2 0 0 0 0 13 27 0 0 2
465 232
465 225
1 0 0 0 0 0 0 23 0 0 16 2
550 212
517 212
5 1 0 0 0 0 0 27 24 0 0 3
483 212
517 212
517 206
0 1 0 0 0 0 0 0 27 19 0 2
409 206
447 206
1 4 0 0 0 0 0 32 27 0 0 2
465 178
465 199
5 0 0 0 0 0 0 26 0 0 20 3
272 245
409 245
409 205
1 1 0 0 0 0 0 39 20 0 0 3
346 205
414 205
414 201
1 2 0 0 0 0 0 22 39 0 0 3
313 133
313 205
326 205
1 2 0 0 0 0 0 30 20 0 0 2
414 160
414 165
1 0 0 0 0 0 0 22 0 0 24 2
313 133
313 133
5 1 0 0 0 0 0 25 21 0 0 2
277 133
338 133
1 2 0 0 0 0 0 26 19 0 0 2
236 251
236 314
0 0 0 0 0 0 0 0 0 30 46 3
109 213
109 214
224 214
2 2 0 0 0 0 0 25 16 0 0 3
241 127
181 127
181 314
2 1 0 0 0 0 0 19 18 0 0 4
236 314
249 314
249 315
245 315
2 1 0 0 0 0 0 16 19 0 0 2
181 314
200 314
0 0 0 0 0 0 0 0 0 32 31 3
73 211
73 213
109 213
1 2 0 0 0 0 0 37 38 0 0 2
109 187
109 241
2 0 0 0 0 0 0 15 0 0 33 2
62 211
73 211
1 2 0 0 0 0 0 17 14 0 0 2
73 190
73 232
1 1 0 0 0 0 0 46 45 0 0 2
655 194
613 194
1 3 7 0 0 0 0 33 45 0 0 2
613 139
613 158
2 2 8 0 0 0 0 45 23 0 0 3
590 176
590 212
586 212
1 2 10 0 0 0 0 29 24 0 0 2
517 164
517 170
2 2 14 0 0 0 0 21 1 0 0 4
374 133
456 133
456 71
591 71
1 2 18 0 0 0 0 31 22 0 0 2
313 65
313 97
1 2 21 0 0 0 0 35 18 0 0 2
306 315
281 315
1 1 2 0 0 0 0 16 42 0 0 3
145 314
140 314
140 320
1 3 22 0 0 0 0 34 26 0 0 2
254 225
254 232
1 4 2 0 0 0 0 44 26 0 0 4
254 262
254 267
254 267
254 258
1 4 2 0 0 0 0 41 25 0 0 2
259 152
259 146
1 3 23 0 0 0 0 36 25 0 0 4
259 107
259 106
259 106
259 120
1 2 24 0 0 0 0 25 26 0 0 4
241 139
224 139
224 239
236 239
1 0 2 0 0 0 0 43 0 0 48 3
30 293
30 288
93 288
1 1 2 0 0 0 0 14 38 0 0 6
73 268
73 288
93 288
93 289
109 289
109 261
2 0 25 0 0 0 0 37 0 0 50 3
109 167
109 128
93 128
1 2 25 0 0 0 0 28 17 0 0 4
93 97
93 128
73 128
73 154
1 1 3 0 0 0 0 15 40 0 0 4
26 211
24 211
24 211
26 211
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
255 198 280 222
263 206 271 222
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
259 78 288 102
269 86 277 102
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
450 268 479 292
460 276 468 292
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
257 255 294 279
267 263 283 279
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
264 146 301 170
274 154 290 170
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
460 344 497 368
470 352 486 368
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
468 225 505 249
478 233 494 249
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
418 290 455 314
428 298 444 314
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
415 320 452 344
425 328 441 344
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
434 181 463 205
444 189 452 205
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
433 213 462 237
443 221 451 237
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
217 245 246 269
227 253 235 269
1 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
222 214 251 238
232 222 240 238
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
460 152 489 176
470 160 478 176
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
228 132 257 156
238 140 246 156
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
227 102 256 126
237 110 245 126
1 4
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
