CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 265 204 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89821e-315 0
0
2 +V
167 359 428 0 1 3
0 7
0
0 0 53360 90
3 10V
6 -2 27 6
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.89821e-315 5.26354e-315
0
7 Ground~
168 492 425 0 1 3
0 2
0
0 0 53360 90
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89821e-315 5.30499e-315
0
12 SPST Switch~
165 440 426 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
5 reset
-34 5 1 13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3421 0 0
2
5.89821e-315 5.32571e-315
0
5 4071~
219 414 356 0 3 22
0 8 2 9
0
0 0 112 90
4 4071
-7 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
8157 0 0
2
5.89821e-315 5.34643e-315
0
5 4081~
219 369 381 0 3 22
0 4 5 8
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
5572 0 0
2
5.89821e-315 5.3568e-315
0
7 Pulser~
4 245 278 0 10 12
0 35 36 10 37 0 0 5 5 6
7
0
0 0 5168 0
0
3 V10
-11 -28 10 -20
15 automatic clock
-52 -28 53 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.89821e-315 5.36716e-315
0
7 Ground~
168 446 290 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
43036.5 0
0
7 Ground~
168 385 287 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
43036.5 1
0
7 Ground~
168 173 289 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
43036.5 2
0
7 Ground~
168 113 295 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
43036.5 3
0
2 +V
167 96 308 0 1 3
0 3
0
0 0 53360 180
3 10V
6 -2 27 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
43036.5 4
0
9 CC 7-Seg~
183 123 51 0 17 19
10 34 33 32 28 31 30 29 38 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3536 0 0
2
5.89821e-315 5.37752e-315
0
7 Ground~
168 132 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89821e-315 5.38788e-315
0
2 +V
167 418 202 0 1 3
0 13
0
0 0 53360 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
5.89821e-315 5.39306e-315
0
2 +V
167 141 202 0 1 3
0 14
0
0 0 53360 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89821e-315 5.39824e-315
0
7 Ground~
168 409 205 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.89821e-315 5.40342e-315
0
9 CC 7-Seg~
183 400 53 0 17 19
10 24 23 22 18 21 20 19 39 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9323 0 0
2
5.89821e-315 5.4086e-315
0
4 4511
219 400 157 0 20 29
0 4 17 16 15 2 13 12 19 20
21 18 22 23 24 0 0 0 0 0
6
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
317 0 0
2
5.89821e-315 5.41378e-315
0
4 4029
219 411 245 0 20 29
0 2 2 2 2 9 10 2 2 2
11 15 16 17 4 0 0 0 0 0
6
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
3108 0 0
2
5.89821e-315 5.41896e-315
0
7 Ground~
168 358 36 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4299 0 0
2
5.89821e-315 5.42414e-315
0
7 Ground~
168 164 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
5.89821e-315 5.42933e-315
0
4 4029
219 134 246 0 20 29
0 3 2 2 2 9 10 11 2 2
40 25 26 27 5 0 0 0 0 0
6
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
43036.5 5
0
4 4511
219 123 158 0 20 29
0 5 27 26 25 2 14 12 29 30
31 28 32 33 34 0 0 0 0 0
6
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
43036.5 6
0
13 SemiResistor~
219 397 426 0 4 5
0 2 7 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R6
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
5.89821e-315 5.43192e-315
0
55
3 1 2 0 0 8192 0 23 11 0 0 3
114 280
113 280
113 289
3 4 2 0 0 0 0 23 23 0 0 2
114 280
123 280
2 3 2 0 0 0 0 23 23 0 0 2
105 280
114 280
1 1 3 0 0 4224 0 23 12 0 0 2
96 280
96 293
0 1 4 0 0 8320 0 0 6 36 0 4
373 195
332 195
332 372
345 372
0 2 5 0 0 12416 0 0 6 48 0 4
96 194
68 194
68 390
345 390
2 2 2 0 0 4224 6 5 4 0 0 3
426 372
426 426
423 426
1 1 2 0 0 4096 0 3 4 0 0 2
485 426
457 426
2 1 2 0 0 0 6 4 25 0 0 2
423 426
415 426
2 1 7 0 0 4224 0 25 2 0 0 2
379 426
370 426
3 1 8 0 0 4224 0 6 5 0 0 3
390 381
408 381
408 372
3 0 9 0 0 4096 0 5 0 0 14 2
417 326
417 327
3 0 10 0 0 8192 0 7 0 0 20 3
269 269
289 269
289 314
5 5 9 0 0 8320 0 23 20 0 0 4
141 280
141 327
418 327
418 279
9 1 2 0 0 0 0 23 10 0 0 3
177 280
177 283
173 283
8 1 2 0 0 0 0 23 10 0 0 3
168 280
168 283
173 283
9 1 2 0 0 0 0 20 8 0 0 3
454 279
454 284
446 284
8 1 2 0 0 0 0 20 8 0 0 3
445 279
445 284
446 284
7 1 2 0 0 0 0 20 8 0 0 3
436 285
436 284
446 284
6 6 10 0 0 8320 0 23 20 0 0 4
150 280
150 314
427 314
427 279
7 10 11 0 0 8320 0 23 20 0 0 5
159 286
159 303
471 303
471 209
418 209
1 0 2 0 0 0 0 9 0 0 24 3
385 281
385 279
386 279
4 3 2 0 0 0 0 20 20 0 0 2
400 279
391 279
3 2 2 0 0 0 0 20 20 0 0 2
391 279
382 279
1 2 2 0 0 0 0 20 20 0 0 2
373 279
382 279
1 0 12 0 0 12288 0 1 0 0 27 6
266 191
266 192
266 192
266 180
265 180
265 181
7 7 12 0 0 4224 0 24 19 0 0 3
150 181
427 181
427 180
6 1 13 0 0 4224 0 19 15 0 0 4
418 180
418 188
418 188
418 187
5 1 2 0 0 0 0 19 17 0 0 2
409 180
409 199
6 1 14 0 0 4224 0 24 16 0 0 4
141 181
141 189
141 189
141 187
5 1 2 0 0 0 0 24 14 0 0 2
132 181
132 197
9 1 2 0 0 8320 0 18 21 0 0 4
400 11
400 7
358 7
358 30
4 11 15 0 0 4224 0 19 20 0 0 2
400 174
400 215
3 12 16 0 0 4224 0 19 20 0 0 2
391 174
391 215
2 13 17 0 0 4224 0 19 20 0 0 2
382 174
382 215
1 14 4 0 0 0 0 19 20 0 0 2
373 174
373 215
4 11 18 0 0 4224 0 18 19 0 0 3
397 89
397 110
400 110
7 8 19 0 0 4224 0 18 19 0 0 4
415 89
415 103
427 103
427 110
6 9 20 0 0 4224 0 18 19 0 0 4
409 89
409 108
418 108
418 110
5 10 21 0 0 4224 0 18 19 0 0 3
403 89
403 110
409 110
3 12 22 0 0 4224 0 18 19 0 0 2
391 89
391 110
2 13 23 0 0 4224 0 18 19 0 0 3
385 89
385 110
382 110
1 14 24 0 0 4224 0 18 19 0 0 3
379 89
379 110
373 110
9 1 2 0 0 0 0 13 22 0 0 4
123 9
123 6
164 6
164 22
4 11 25 0 0 4224 0 24 23 0 0 2
123 175
123 216
3 12 26 0 0 4224 0 24 23 0 0 2
114 175
114 216
2 13 27 0 0 4224 0 24 23 0 0 2
105 175
105 216
1 14 5 0 0 0 0 24 23 0 0 2
96 175
96 216
4 11 28 0 0 4224 0 13 24 0 0 4
120 87
120 112
123 112
123 111
7 8 29 0 0 4224 0 13 24 0 0 4
138 87
138 102
150 102
150 111
6 9 30 0 0 4224 0 13 24 0 0 4
132 87
132 107
141 107
141 111
5 10 31 0 0 4224 0 13 24 0 0 4
126 87
126 112
132 112
132 111
3 12 32 0 0 4224 0 13 24 0 0 2
114 87
114 111
2 13 33 0 0 4224 0 13 24 0 0 4
108 87
108 112
105 112
105 111
1 14 34 0 0 4224 0 13 24 0 0 4
102 87
102 112
96 112
96 111
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
