CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 80 10
176 79 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 166 111 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 U2
-13 -21 1 -13
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89827e-315 0
0
13 Logic Switch~
5 41 303 0 1 11
0 12
0
0 0 21088 0
2 0V
-6 -16 8 -8
2 U1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89827e-315 0
0
2 +V
167 1062 306 0 1 3
0 7
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89827e-315 0
0
14 NO PushButton~
191 1095 371 0 2 5
0 35 7
0
0 0 4704 0
0
2 U1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 512 1 0 0 0
1 S
3421 0 0
2
5.89827e-315 0
0
14 NO PushButton~
191 1178 151 0 2 5
0 36 8
0
0 0 4704 0
0
3 U12
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 512 1 0 0 0
1 S
8157 0 0
2
5.89827e-315 5.26354e-315
0
2 +V
167 1107 104 0 1 3
0 8
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
5.89827e-315 0
0
5 4011~
219 283 132 0 3 22
0 5 6 4
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 9 0
1 U
8901 0 0
2
5.89827e-315 0
0
5 4011~
219 270 53 0 3 22
0 10 4 5
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 9 0
1 U
7361 0 0
2
5.89827e-315 5.30499e-315
0
14 NO PushButton~
191 1257 385 0 2 5
0 37 11
0
0 0 4704 0
0
2 U2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 512 1 0 0 0
1 S
4747 0 0
2
5.89827e-315 5.26354e-315
0
2 +V
167 1229 337 0 1 3
0 11
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.89827e-315 0
0
5 4011~
219 188 332 0 3 22
0 9 12 3
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 9 0
1 U
3472 0 0
2
43108.6 0
0
5 4011~
219 171 233 0 3 22
0 10 3 9
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 9 0
1 U
9998 0 0
2
43108.6 1
0
7 Ground~
168 357 740 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
43108.6 2
0
7 Ground~
168 324 742 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
43108.6 3
0
5 4073~
219 582 350 0 4 22
0 14 28 27 23
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
3835 0 0
2
5.89827e-315 5.30499e-315
0
5 4073~
219 582 285 0 4 22
0 14 15 5 31
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
3670 0 0
2
5.89827e-315 5.32571e-315
0
5 4073~
219 582 386 0 4 22
0 26 25 5 20
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
5616 0 0
2
5.89827e-315 5.34643e-315
0
5 4073~
219 582 420 0 4 22
0 14 5 9 21
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
9323 0 0
2
5.89827e-315 5.3568e-315
0
12 D Flip-Flop~
219 601 581 0 4 9
0 19 10 38 13
0
0 0 5216 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
12 F.F. D (X 1)
-44 -68 40 -60
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
5.89827e-315 5.36716e-315
0
12 D Flip-Flop~
219 488 583 0 4 9
0 18 10 39 14
0
0 0 5216 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
12 F.F. D (X 2)
-39 -56 45 -48
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
5.89827e-315 5.37752e-315
0
5 4071~
219 788 535 0 3 22
0 14 13 17
0
0 0 1120 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
1 Y
33 -21 40 -13
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
4299 0 0
2
5.89827e-315 5.38788e-315
0
8 4-In OR~
219 665 400 0 5 22
0 23 20 21 22 18
0
0 0 1120 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
7 X2(t+1)
-13 -26 36 -18
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
9672 0 0
2
5.89827e-315 5.39306e-315
0
5 4049~
219 509 455 0 2 22
0 5 24
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
3 X 2
-88 -79 -67 -71
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
7876 0 0
2
5.89827e-315 5.39824e-315
0
5 4049~
219 499 160 0 2 22
0 14 34
0
0 0 1120 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
3 X 2
-125 -44 -104 -36
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
6369 0 0
2
5.89827e-315 5.40342e-315
0
5 4049~
219 476 377 0 2 22
0 13 26
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
3 X 1
-91 -146 -70 -138
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
9172 0 0
2
5.89827e-315 5.4086e-315
0
5 4049~
219 473 350 0 2 22
0 9 28
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
7100 0 0
2
5.89827e-315 5.41378e-315
0
5 4049~
219 500 217 0 2 22
0 9 33
0
0 0 1120 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
3 X 1
-100 -102 -79 -94
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 4 0
1 U
3820 0 0
2
5.89827e-315 5.41896e-315
0
5 4049~
219 511 359 0 2 22
0 5 27
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
7678 0 0
2
5.89827e-315 5.42414e-315
0
5 4081~
219 582 208 0 3 22
0 13 33 29
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
3 X 1
-339 -134 -318 -126
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
5.89827e-315 5.42933e-315
0
5 4081~
219 582 248 0 3 22
0 13 5 30
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
3 U 2
-374 -90 -353 -82
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3178 0 0
2
5.89827e-315 5.43192e-315
0
5 4073~
219 581 169 0 4 22
0 34 13 40 32
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 1 2 0
1 U
3409 0 0
2
5.89827e-315 5.43451e-315
0
5 4073~
219 582 455 0 4 22
0 13 24 9 22
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
3 U 1
-413 -51 -392 -43
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 70
65 0 0 0 3 1 1 0
1 U
3951 0 0
2
5.89827e-315 5.4371e-315
0
8 4-In OR~
219 666 225 0 5 22
0 32 29 30 31 19
0
0 0 1120 0
4 4072
-14 -24 14 -16
3 U9B
-3 -25 18 -17
7 X1(t+1)
-11 -26 38 -18
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
8885 0 0
2
5.89827e-315 5.43969e-315
0
5 4049~
219 512 386 0 2 22
0 9 25
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
3 X 1
-91 -146 -70 -138
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
3780 0 0
2
5.89827e-315 5.44228e-315
0
4 LED~
171 860 534 0 2 2
12 17 2
0
0 0 96 90
4 LED1
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9265 0 0
2
5.89827e-315 5.44487e-315
0
7 Ground~
168 892 555 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9442 0 0
2
5.89827e-315 5.44746e-315
0
4 LED~
171 845 454 0 2 2
10 16 17
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9424 0 0
2
5.89827e-315 5.45005e-315
0
2 +V
167 845 390 0 1 3
0 16
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9968 0 0
2
5.89827e-315 5.45264e-315
0
5 4069~
219 484 285 0 2 22
0 9 15
0
0 0 608 0
4 4069
-7 -24 21 -16
4 U10A
-14 -20 14 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
9281 0 0
2
5.89827e-315 5.45523e-315
0
7 Pulser~
4 68 562 0 10 12
0 41 42 10 43 0 0 10 10 9
8
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8464 0 0
2
5.89827e-315 5.45782e-315
0
9 Resistor~
219 357 699 0 3 5
0 2 5 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
43108.6 4
0
9 Resistor~
219 329 697 0 3 5
0 2 9 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
43108.6 5
0
70
3 2 3 0 0 8320 0 11 12 0 0 5
215 332
215 279
84 279
84 242
147 242
0 2 4 0 0 4096 0 0 8 3 0 4
209 69
238 69
238 62
246 62
3 0 4 0 0 8320 0 7 0 0 0 4
310 132
310 102
209 102
209 65
0 0 5 0 0 4096 0 0 0 10 68 2
297 76
326 76
1 0 6 0 0 8192 0 1 0 0 12 4
178 111
192 111
192 137
191 137
1 2 7 0 0 8320 0 3 4 0 0 4
1062 315
1061 315
1061 379
1078 379
1 2 8 0 0 8320 0 6 5 0 0 3
1107 113
1107 159
1161 159
0 0 9 0 0 4096 0 0 0 18 9 3
211 260
302 260
302 206
2 0 9 0 0 8320 0 42 0 0 0 4
329 679
321 679
321 206
292 206
1 3 5 0 0 4096 0 7 8 0 0 4
259 123
259 84
297 84
297 53
1 0 10 0 0 8192 0 8 0 0 14 4
246 44
228 44
228 387
117 387
0 2 6 0 0 8320 0 0 7 0 0 4
191 141
191 133
259 133
259 141
1 2 11 0 0 4224 0 10 9 0 0 3
1229 346
1229 393
1240 393
1 0 10 0 0 0 0 12 0 0 16 3
147 224
117 224
117 565
1 2 12 0 0 4224 0 2 11 0 0 5
53 303
126 303
126 297
164 297
164 341
2 3 10 0 0 4224 0 20 40 0 0 4
464 565
106 565
106 553
92 553
0 2 10 0 0 0 0 0 19 16 0 4
434 565
434 582
577 582
577 563
3 1 9 0 0 0 0 12 11 0 0 8
198 233
200 233
200 247
211 247
211 263
111 263
111 323
164 323
1 1 2 0 0 4096 0 13 41 0 0 2
357 734
357 717
1 1 2 0 0 4224 0 14 42 0 0 3
324 736
324 715
329 715
4 0 13 0 0 12288 0 19 0 0 70 4
625 545
655 545
655 500
409 500
4 0 14 0 0 12288 0 20 0 0 69 4
512 547
534 547
534 516
387 516
1 0 14 0 0 12288 0 21 0 0 69 4
775 526
742 526
742 484
387 484
2 0 13 0 0 12288 0 21 0 0 70 4
775 544
750 544
750 635
409 635
1 0 9 0 0 0 0 39 0 0 9 4
469 285
344 285
344 286
321 286
2 2 15 0 0 4224 0 39 16 0 0 2
505 285
558 285
1 0 13 0 0 0 0 30 0 0 70 2
558 239
409 239
1 1 16 0 0 4224 0 38 37 0 0 2
845 399
845 444
0 2 17 0 0 4224 0 0 37 31 0 2
845 535
845 464
2 1 2 0 0 0 0 35 36 0 0 3
873 535
892 535
892 549
3 1 17 0 0 0 0 21 35 0 0 2
821 535
853 535
5 1 18 0 0 8320 0 22 20 0 0 5
698 400
698 590
455 590
455 547
464 547
5 1 19 0 0 8320 0 33 19 0 0 6
699 225
727 225
727 607
566 607
566 545
577 545
4 2 20 0 0 4224 0 17 22 0 0 4
603 386
634 386
634 396
648 396
4 3 21 0 0 4224 0 18 22 0 0 4
603 420
635 420
635 405
648 405
4 4 22 0 0 4224 0 32 22 0 0 3
603 455
648 455
648 414
4 1 23 0 0 4224 0 15 22 0 0 3
603 350
648 350
648 387
3 0 9 0 0 0 0 32 0 0 9 2
558 464
321 464
1 0 5 0 0 4096 0 23 0 0 68 2
494 455
358 455
2 2 24 0 0 4224 0 32 23 0 0 2
558 455
530 455
1 0 13 0 0 0 0 32 0 0 70 2
558 446
409 446
3 0 9 0 0 0 0 18 0 0 9 2
558 429
321 429
2 0 5 0 0 4096 0 18 0 0 68 2
558 420
358 420
1 0 14 0 0 0 0 18 0 0 69 2
558 411
387 411
3 0 5 0 0 0 0 17 0 0 68 2
558 395
358 395
1 0 9 0 0 0 0 34 0 0 9 2
497 386
321 386
2 2 25 0 0 4224 0 34 17 0 0 2
533 386
558 386
1 0 13 0 0 0 0 25 0 0 70 2
461 377
409 377
1 2 26 0 0 4224 0 17 25 0 0 2
558 377
497 377
1 0 5 0 0 0 0 28 0 0 68 2
496 359
358 359
3 2 27 0 0 4224 0 15 28 0 0 2
558 359
532 359
1 0 9 0 0 0 0 26 0 0 9 2
458 350
321 350
2 2 28 0 0 4224 0 15 26 0 0 2
558 350
494 350
1 0 14 0 0 0 0 15 0 0 69 2
558 341
387 341
3 2 29 0 0 4224 0 29 33 0 0 4
603 208
637 208
637 221
649 221
3 3 30 0 0 4224 0 30 33 0 0 4
603 248
638 248
638 230
649 230
4 4 31 0 0 4224 0 16 33 0 0 3
603 285
649 285
649 239
4 1 32 0 0 4224 0 31 33 0 0 3
602 169
649 169
649 212
3 0 5 0 0 0 0 16 0 0 68 2
558 294
358 294
1 0 14 0 0 0 0 16 0 0 69 2
558 276
387 276
2 0 5 0 0 0 0 30 0 0 68 2
558 257
358 257
2 2 33 0 0 4224 0 27 29 0 0 2
521 217
558 217
1 0 13 0 0 0 0 29 0 0 70 2
558 199
409 199
0 1 9 0 0 0 0 0 27 9 0 2
321 217
485 217
0 2 13 0 0 0 0 0 31 70 0 2
409 169
557 169
2 1 34 0 0 4224 0 24 31 0 0 2
520 160
557 160
0 1 14 0 0 0 0 0 24 69 0 2
387 160
484 160
0 2 5 0 0 28800 0 0 41 0 0 9
326 102
326 27
367 27
367 103
353 103
353 143
358 143
358 681
357 681
0 0 14 0 0 4224 0 0 0 0 0 2
387 137
387 684
0 0 13 0 0 4224 0 0 0 0 0 2
409 137
409 684
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
