CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 18 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
31
6 Diode~
219 149 88 0 2 5
0 19 25
0
0 0 64 90
6 1N4148
12 0 54 8
2 D6
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
5130 0 0
2
5.89839e-315 5.46041e-315
0
7 Ground~
168 83 248 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
5.89839e-315 5.45782e-315
0
7 Ground~
168 179 518 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89839e-315 5.45523e-315
0
7 Ground~
168 31 521 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.89839e-315 5.45264e-315
0
14 NO PushButton~
191 23 484 0 2 5
0 3 2
0
0 0 4192 90
0
2 S1
15 -5 29 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8157 0 0
2
5.89839e-315 5.45005e-315
0
5 7474~
219 276 343 0 6 22
0 5 11 6 10 14 18
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 3 0
1 U
5572 0 0
2
5.89839e-315 5.44746e-315
0
5 7474~
219 389 343 0 6 22
0 8 18 6 5 4 17
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 3 0
1 U
8901 0 0
2
5.89839e-315 5.44487e-315
0
5 7474~
219 499 343 0 6 22
0 5 17 6 9 13 16
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 2 0
1 U
7361 0 0
2
5.89839e-315 5.44228e-315
0
5 7474~
219 601 343 0 6 22
0 7 16 6 5 12 11
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 2 0
1 U
4747 0 0
2
5.89839e-315 5.43969e-315
0
9 Inverter~
13 176 375 0 2 22
0 3 6
0
0 0 96 90
5 74F04
-18 -19 17 -11
3 U1C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
972 0 0
2
5.89839e-315 5.4371e-315
0
9 Inverter~
13 256 154 0 2 22
0 24 5
0
0 0 96 0
5 74F04
-18 -19 17 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3472 0 0
2
5.89839e-315 5.43451e-315
0
9 Inverter~
13 174 154 0 2 22
0 19 24
0
0 0 96 0
5 74F04
-18 -19 17 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9998 0 0
2
5.89839e-315 5.43192e-315
0
4 LED~
171 346 141 0 2 2
10 23 14
0
0 0 112 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3536 0 0
2
5.89839e-315 5.42933e-315
0
4 LED~
171 426 141 0 2 2
10 22 4
0
0 0 112 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4597 0 0
2
5.89839e-315 5.42414e-315
0
4 LED~
171 639 144 0 2 2
10 20 12
0
0 0 112 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3835 0 0
2
5.89839e-315 5.41896e-315
0
4 LED~
171 534 141 0 2 2
10 21 13
0
0 0 112 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3670 0 0
2
5.89839e-315 5.41378e-315
0
2 +V
167 601 233 0 1 3
0 7
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
5.89839e-315 5.4086e-315
0
2 +V
167 499 391 0 1 3
0 9
0
0 0 53472 180
3 10V
-11 -22 10 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
5.89839e-315 5.40342e-315
0
2 +V
167 389 237 0 1 3
0 8
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
5.89839e-315 5.39824e-315
0
2 +V
167 149 29 0 1 3
0 25
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
5.89839e-315 5.39306e-315
0
2 +V
167 83 34 0 1 3
0 26
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.89839e-315 5.38788e-315
0
2 +V
167 31 392 0 1 3
0 15
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
5.89839e-315 5.37752e-315
0
2 +V
167 346 27 0 1 3
0 23
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
5.89839e-315 5.36716e-315
0
2 +V
167 276 395 0 1 3
0 10
0
0 0 53472 180
3 10V
-12 -22 9 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6369 0 0
2
5.89839e-315 5.3568e-315
0
2 +V
167 534 26 0 1 3
0 21
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9172 0 0
2
5.89839e-315 5.34643e-315
0
2 +V
167 639 25 0 1 3
0 20
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
5.89839e-315 5.32571e-315
0
2 +V
167 426 25 0 1 3
0 22
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3820 0 0
2
5.89839e-315 5.30499e-315
0
10 Polar Cap~
219 180 486 0 2 5
0 3 2
0
0 0 64 270
5 10 uF
3 4 38 12
2 C2
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7678 0 0
2
5.89839e-315 5.26354e-315
0
10 Polar Cap~
219 84 191 0 2 5
0 19 2
0
0 0 64 782
5 10 uF
3 4 38 12
2 C1
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
961 0 0
2
5.89839e-315 0
0
9 Resistor~
219 83 89 0 4 5
0 19 26 0 1
0
0 0 96 90
4 56 K
1 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
5.89839e-315 5.46559e-315
0
9 Resistor~
219 31 424 0 4 5
0 3 15 0 1
0
0 0 96 90
4 68 K
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.89839e-315 5.463e-315
0
37
0 0 3 0 0 4224 0 0 0 21 23 2
31 454
179 454
2 5 4 0 0 4224 0 14 7 0 0 3
426 151
426 325
419 325
1 0 5 0 0 4096 0 6 0 0 6 2
276 280
276 208
2 0 5 0 0 0 0 11 0 0 6 3
277 154
334 154
334 208
4 0 5 0 0 0 0 7 0 0 6 2
389 355
389 423
4 1 5 0 0 8320 0 9 8 0 0 6
601 355
601 423
229 423
229 208
499 208
499 280
0 2 6 0 0 4096 0 0 10 10 0 3
248 341
179 341
179 357
3 0 6 0 0 8192 0 8 0 0 10 3
475 325
444 325
444 405
3 0 6 0 0 0 0 7 0 0 10 3
365 325
348 325
348 405
3 3 6 0 0 12416 0 6 9 0 0 6
252 325
248 325
248 405
569 405
569 325
577 325
1 1 7 0 0 4224 0 17 9 0 0 2
601 242
601 280
1 1 8 0 0 4224 0 19 7 0 0 2
389 246
389 280
4 1 9 0 0 4224 0 8 18 0 0 2
499 355
499 376
4 1 10 0 0 4224 0 6 24 0 0 2
276 355
276 380
2 6 11 0 0 12416 0 6 9 0 0 6
252 307
181 307
181 184
721 184
721 307
625 307
2 5 12 0 0 4224 0 15 9 0 0 3
639 154
639 325
631 325
2 5 13 0 0 4224 0 16 8 0 0 3
534 151
534 325
529 325
2 5 14 0 0 4224 0 13 6 0 0 3
346 151
346 325
306 325
1 2 15 0 0 4224 0 22 31 0 0 2
31 401
31 406
2 1 2 0 0 4096 0 5 4 0 0 2
31 501
31 515
1 1 3 0 0 0 0 31 5 0 0 2
31 442
31 467
2 1 2 0 0 4096 0 28 3 0 0 2
179 493
179 512
1 1 3 0 0 0 0 10 28 0 0 2
179 393
179 476
6 2 16 0 0 4224 0 8 9 0 0 2
523 307
577 307
6 2 17 0 0 4224 0 7 8 0 0 2
413 307
475 307
6 2 18 0 0 4224 0 6 7 0 0 2
300 307
365 307
1 0 19 0 0 4096 0 1 0 0 32 4
149 98
149 149
150 149
150 154
1 1 20 0 0 4224 0 26 15 0 0 2
639 34
639 134
1 1 21 0 0 4224 0 25 16 0 0 2
534 35
534 131
1 1 22 0 0 4224 0 27 14 0 0 2
426 34
426 131
1 1 23 0 0 4224 0 23 13 0 0 2
346 36
346 131
0 1 19 0 0 4224 0 0 12 34 0 2
83 154
159 154
2 1 24 0 0 4224 0 12 11 0 0 2
195 154
241 154
1 1 19 0 0 0 0 30 29 0 0 2
83 107
83 181
2 1 2 0 0 4224 0 29 2 0 0 2
83 198
83 242
1 2 25 0 0 4224 0 20 1 0 0 2
149 38
149 78
1 2 26 0 0 4224 0 21 30 0 0 2
83 43
83 71
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
