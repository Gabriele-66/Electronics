CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 120 10
176 80 1313 661
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 675 194 0 1 11
0 6
0
0 0 20592 270
2 0V
11 0 25 8
2 V2
11 -10 25 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89821e-315 0
0
13 Logic Switch~
5 265 204 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
9 lamp test
-29 15 34 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89821e-315 0
0
7 Pulser~
4 245 272 0 10 12
0 40 41 3 42 0 0 5 5 1
7
0
0 0 5168 0
0
3 V10
-11 -28 10 -20
15 automatic clock
-52 -28 53 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9281 0 0
2
43033.9 0
0
2 +V
167 556 100 0 1 3
0 4
0
0 0 53360 90
3 10V
6 -2 27 6
2 V1
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
43033.9 2
0
7 Ground~
168 661 97 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
43033.9 1
0
12 SPST Switch~
165 637 98 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
5 clock
-40 -15 -5 -7
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3171 0 0
2
43033.9 0
0
2 +V
167 338 434 0 1 3
0 8
0
0 0 53360 90
3 10V
6 -2 27 6
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89821e-315 5.30499e-315
0
7 Ground~
168 471 431 0 1 3
0 2
0
0 0 53360 90
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
5.89821e-315 5.26354e-315
0
12 SPST Switch~
165 419 432 0 10 11
0 2 2 0 0 0 0 0 0 0
1
0
0 0 4720 0
0
6 preset
-37 5 5 13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5283 0 0
2
5.89821e-315 0
0
5 4071~
219 393 361 0 3 22
0 11 2 12
0
0 0 112 90
4 4071
-7 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
6874 0 0
2
5.89821e-315 0
0
9 4-In NOR~
219 314 245 0 5 22
0 16 15 14 13 10
0
0 0 112 270
4 4002
-14 -24 14 -16
3 U7B
29 -8 50 0
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 4 0
1 U
5305 0 0
2
5.89821e-315 0
0
9 4-In NOR~
219 48 238 0 5 22
0 20 19 18 17 9
0
0 0 112 270
4 4002
-14 -24 14 -16
3 U7A
29 -8 50 0
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 4 0
1 U
34 0 0
2
5.89821e-315 0
0
5 4081~
219 366 391 0 3 22
0 10 9 11
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
969 0 0
2
5.89821e-315 5.37752e-315
0
5 4011~
219 736 44 0 3 22
0 43 44 45
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 512 4 1 3 0
1 U
8402 0 0
2
5.89821e-315 5.36716e-315
0
5 4001~
219 639 320 0 3 22
0 46 47 48
0
0 0 624 270
4 4001
-14 -24 14 -16
3 U9A
31 -10 52 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 512 4 1 6 0
1 U
3751 0 0
2
5.89821e-315 0
0
5 4011~
219 824 335 0 3 22
0 49 50 51
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U5B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 512 4 2 3 0
1 U
4292 0 0
2
5.89821e-315 0
0
8 4-In OR~
219 733 328 0 5 22
0 52 53 54 55 56
0
0 0 624 270
4 4072
-14 -24 14 -16
3 U8A
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 5 0
1 U
6118 0 0
2
5.89821e-315 0
0
7 Ground~
168 446 290 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
34 0 0
2
43033.9 0
0
7 Ground~
168 385 287 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
43033.9 1
0
7 Ground~
168 173 289 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
319 0 0
2
43033.9 2
0
7 Ground~
168 96 307 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3976 0 0
2
43033.9 3
0
2 +V
167 109 299 0 1 3
0 22
0
0 0 53360 180
3 10V
6 -2 27 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7634 0 0
2
43033.9 4
0
9 CC 7-Seg~
183 123 51 0 17 19
10 39 38 37 33 36 35 34 57 2
0 1 1 0 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
523 0 0
2
5.89821e-315 5.26354e-315
0
7 Ground~
168 132 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6748 0 0
2
5.89821e-315 5.30499e-315
0
2 +V
167 418 202 0 1 3
0 24
0
0 0 53360 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6901 0 0
2
5.89821e-315 5.32571e-315
0
2 +V
167 141 202 0 1 3
0 25
0
0 0 53360 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
842 0 0
2
5.89821e-315 5.34643e-315
0
7 Ground~
168 409 205 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3277 0 0
2
5.89821e-315 5.3568e-315
0
9 CC 7-Seg~
183 400 53 0 17 19
10 32 31 30 26 29 28 27 58 2
0 0 1 1 1 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4212 0 0
2
5.89821e-315 5.36716e-315
0
4 4511
219 400 157 0 20 29
0 16 15 14 13 2 24 23 27 28
29 26 30 31 32 0 0 0 0 0
6
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4720 0 0
2
5.89821e-315 5.37752e-315
0
4 4029
219 411 245 0 20 29
0 2 2 2 2 12 3 2 2 2
21 13 14 15 16 0 0 0 0 0
6
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
5551 0 0
2
5.89821e-315 5.38788e-315
0
7 Ground~
168 358 36 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
5.89821e-315 5.39306e-315
0
7 Ground~
168 164 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8745 0 0
2
5.89821e-315 5.39824e-315
0
4 4029
219 134 246 0 20 29
0 2 22 22 2 12 3 21 2 2
59 17 18 19 20 0 0 0 0 0
4
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 512 1 0 0 0
1 U
9592 0 0
2
43033.9 5
0
4 4511
219 123 158 0 20 29
0 20 19 18 17 2 25 23 34 35
36 33 37 38 39 0 0 0 0 0
4
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8748 0 0
2
43033.9 6
0
13 SemiResistor~
219 594 98 0 4 5
0 2 4 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R5
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
43033.9 3
0
13 SemiResistor~
219 376 432 0 4 5
0 2 8 0 1
0
0 0 80 180
8 RESISTOR
8 0 64 8
2 R6
29 -10 43 -2
0
0
14 %D %1 %2 %M 1K
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
5.89821e-315 5.32571e-315
0
68
3 0 3 0 0 8208 0 3 0 0 29 3
269 263
290 263
290 314
1 2 4 0 0 4224 0 4 35 0 0 2
567 98
576 98
0 0 2 0 0 4224 5 0 0 0 5 2
615 149
615 98
1 1 2 0 0 4096 0 5 6 0 0 4
654 98
660 98
660 98
654 98
2 1 2 0 0 0 5 6 35 0 0 2
620 98
612 98
0 1 6 0 0 8320 0 0 1 0 0 3
676 231
675 231
675 206
2 2 2 0 0 4224 7 10 9 0 0 3
405 377
405 432
402 432
1 1 2 0 0 4096 0 8 9 0 0 2
464 432
436 432
2 1 2 0 0 0 7 9 36 0 0 2
402 432
394 432
2 1 8 0 0 4224 0 36 7 0 0 2
358 432
349 432
5 2 9 0 0 8320 0 12 13 0 0 3
54 271
54 400
342 400
5 1 10 0 0 4224 0 11 13 0 0 3
320 278
320 382
342 382
1 3 11 0 0 4224 0 10 13 0 0 2
387 377
387 391
0 3 12 0 0 4096 0 0 10 23 0 2
396 327
396 331
4 0 13 0 0 8320 0 11 0 0 46 3
306 222
306 195
400 195
3 0 14 0 0 8320 0 11 0 0 47 3
315 222
315 203
391 203
2 0 15 0 0 8320 0 11 0 0 48 3
324 222
324 210
382 210
1 14 16 0 0 8192 0 11 30 0 0 4
333 222
333 213
373 213
373 215
4 0 17 0 0 8320 0 12 0 0 58 3
40 215
40 191
123 191
3 0 18 0 0 8320 0 12 0 0 59 3
49 215
49 198
114 198
2 0 19 0 0 8320 0 12 0 0 60 3
58 215
58 204
105 204
1 0 20 0 0 8192 0 12 0 0 61 3
67 215
67 211
96 211
5 5 12 0 0 8320 0 33 30 0 0 4
141 280
141 327
418 327
418 279
9 1 2 0 0 0 0 33 20 0 0 3
177 280
177 283
173 283
8 1 2 0 0 0 0 33 20 0 0 3
168 280
168 283
173 283
9 1 2 0 0 0 0 30 18 0 0 3
454 279
454 284
446 284
8 1 2 0 0 0 0 30 18 0 0 3
445 279
445 284
446 284
7 1 2 0 0 0 0 30 18 0 0 3
436 285
436 284
446 284
6 6 3 0 0 8320 0 33 30 0 0 4
150 280
150 314
427 314
427 279
7 10 21 0 0 8320 0 33 30 0 0 5
159 286
159 303
471 303
471 209
418 209
1 4 2 0 0 0 0 21 33 0 0 3
96 301
123 301
123 280
1 1 2 0 0 0 0 33 21 0 0 2
96 280
96 301
1 0 22 0 0 4096 0 22 0 0 34 2
109 284
109 280
2 3 22 0 0 4224 0 33 33 0 0 2
105 280
114 280
1 0 2 0 0 0 0 19 0 0 37 3
385 281
385 279
386 279
4 3 2 0 0 0 0 30 30 0 0 2
400 279
391 279
3 2 2 0 0 0 0 30 30 0 0 2
391 279
382 279
1 2 2 0 0 0 0 30 30 0 0 2
373 279
382 279
1 0 23 0 0 12288 0 2 0 0 40 6
266 191
266 192
266 192
266 180
265 180
265 181
7 7 23 0 0 4224 0 34 29 0 0 3
150 181
427 181
427 180
6 1 24 0 0 4224 0 29 25 0 0 4
418 180
418 188
418 188
418 187
5 1 2 0 0 0 0 29 27 0 0 2
409 180
409 199
6 1 25 0 0 4224 0 34 26 0 0 4
141 181
141 189
141 189
141 187
5 1 2 0 0 0 0 34 24 0 0 2
132 181
132 197
9 1 2 0 0 8320 0 28 31 0 0 4
400 11
400 7
358 7
358 30
4 11 13 0 0 0 0 29 30 0 0 2
400 174
400 215
3 12 14 0 0 0 0 29 30 0 0 2
391 174
391 215
2 13 15 0 0 0 0 29 30 0 0 2
382 174
382 215
1 14 16 0 0 4224 0 29 30 0 0 2
373 174
373 215
4 11 26 0 0 4224 0 28 29 0 0 3
397 89
397 110
400 110
7 8 27 0 0 4224 0 28 29 0 0 4
415 89
415 103
427 103
427 110
6 9 28 0 0 4224 0 28 29 0 0 4
409 89
409 108
418 108
418 110
5 10 29 0 0 4224 0 28 29 0 0 3
403 89
403 110
409 110
3 12 30 0 0 4224 0 28 29 0 0 2
391 89
391 110
2 13 31 0 0 4224 0 28 29 0 0 3
385 89
385 110
382 110
1 14 32 0 0 4224 0 28 29 0 0 3
379 89
379 110
373 110
9 1 2 0 0 0 0 23 32 0 0 4
123 9
123 6
164 6
164 22
4 11 17 0 0 0 0 34 33 0 0 2
123 175
123 216
3 12 18 0 0 0 0 34 33 0 0 2
114 175
114 216
2 13 19 0 0 0 0 34 33 0 0 2
105 175
105 216
1 14 20 0 0 4224 0 34 33 0 0 2
96 175
96 216
4 11 33 0 0 4224 0 23 34 0 0 4
120 87
120 112
123 112
123 111
7 8 34 0 0 4224 0 23 34 0 0 4
138 87
138 102
150 102
150 111
6 9 35 0 0 4224 0 23 34 0 0 4
132 87
132 107
141 107
141 111
5 10 36 0 0 4224 0 23 34 0 0 4
126 87
126 112
132 112
132 111
3 12 37 0 0 4224 0 23 34 0 0 2
114 87
114 111
2 13 38 0 0 4224 0 23 34 0 0 4
108 87
108 112
105 112
105 111
1 14 39 0 0 4224 0 23 34 0 0 4
102 87
102 112
96 112
96 111
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
