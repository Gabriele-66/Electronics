CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 170 30 100 10
176 80 1325 608
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 68 27 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21744 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
3 U 2
-10 -26 11 -18
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
43072.7 0
0
13 Logic Switch~
5 39 27 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
3 U 1
-10 -25 11 -17
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
43072.7 1
0
7 Pulser~
4 204 541 0 10 12
0 26 27 3 28 0 0 5 5 6
7
0
0 0 4656 90
0
2 V3
23 -5 37 3
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7678 0 0
2
43072.8 0
0
7 Ground~
168 602 451 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
961 0 0
2
43072.8 0
0
4 LED~
171 570 430 0 2 2
10 4 2
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3178 0 0
2
43072.8 0
0
5 4049~
219 222 282 0 2 22
0 13 16
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
3 X 1
-91 -146 -70 -138
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
3409 0 0
2
43072.7 0
0
8 4-In OR~
219 376 121 0 5 22
0 23 20 21 22 8
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U9B
-3 -25 18 -17
7 X1(t+1)
-11 -26 38 -18
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
3951 0 0
2
43072.7 4
0
5 4073~
219 292 351 0 4 22
0 5 15 13 11
0
0 0 1136 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
3 U 1
-413 -51 -392 -43
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
8885 0 0
2
43072.7 5
0
5 4073~
219 291 65 0 4 22
0 25 5 13 23
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3780 0 0
2
43072.7 6
0
5 4081~
219 292 144 0 3 22
0 5 14 21
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
3 U 2
-374 -90 -353 -82
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9265 0 0
2
43072.7 7
0
5 4081~
219 292 104 0 3 22
0 5 24 20
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
3 X 1
-339 -134 -318 -126
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9442 0 0
2
43072.7 8
0
5 4049~
219 221 255 0 2 22
0 14 18
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
9424 0 0
2
43072.7 9
0
5 4049~
219 210 113 0 2 22
0 13 24
0
0 0 1136 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
3 X 1
-100 -102 -79 -94
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 4 0
1 U
9968 0 0
2
43072.7 10
0
5 4049~
219 183 246 0 2 22
0 13 19
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
9281 0 0
2
43072.7 11
0
5 4049~
219 186 273 0 2 22
0 5 17
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
3 X 1
-91 -146 -70 -138
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
8464 0 0
2
43072.7 12
0
5 4049~
219 209 56 0 2 22
0 6 25
0
0 0 1136 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
3 X 2
-125 -44 -104 -36
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
7168 0 0
2
43072.7 13
0
5 4049~
219 219 351 0 2 22
0 14 15
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
3 X 2
-88 -79 -67 -71
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
3171 0 0
2
43072.7 15
0
8 4-In OR~
219 375 296 0 5 22
0 12 9 10 11 7
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
7 X2(t+1)
-13 -26 36 -18
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
4139 0 0
2
43072.7 16
0
5 4071~
219 498 431 0 3 22
0 6 5 4
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
1 Y
33 -21 40 -13
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
6435 0 0
2
43072.7 17
0
12 D Flip-Flop~
219 198 479 0 4 9
0 7 3 29 6
0
0 0 5232 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
12 F.F. D (X 2)
-39 -56 45 -48
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5283 0 0
2
43072.7 18
0
12 D Flip-Flop~
219 311 477 0 4 9
0 8 3 30 5
0
0 0 5232 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
12 F.F. D (X 1)
-44 -68 40 -60
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6874 0 0
2
43072.7 19
0
5 4073~
219 292 316 0 4 22
0 6 14 13 10
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
5305 0 0
2
43072.7 20
0
5 4073~
219 292 282 0 4 22
0 17 16 14 9
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
34 0 0
2
43072.7 21
0
5 4073~
219 292 181 0 4 22
0 6 13 14 22
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
969 0 0
2
43072.7 22
0
5 4073~
219 292 246 0 4 22
0 6 19 18 12
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
8402 0 0
2
43072.7 23
0
51
0 2 3 0 0 4224 0 0 21 2 0 4
174 478
254 478
254 459
287 459
2 3 3 0 0 0 0 20 3 0 0 3
174 461
174 517
195 517
2 1 2 0 0 4224 0 5 4 0 0 3
583 431
602 431
602 445
3 1 4 0 0 4224 0 19 5 0 0 2
531 431
563 431
2 0 5 0 0 4096 0 19 0 0 7 2
485 440
355 440
1 0 6 0 0 4096 0 19 0 0 8 2
485 422
246 422
0 4 5 0 0 4096 0 0 21 51 0 4
119 395
355 395
355 441
335 441
0 4 6 0 0 0 0 0 20 50 0 4
97 408
246 408
246 443
222 443
5 1 7 0 0 8320 0 18 20 0 0 5
408 296
408 486
165 486
165 443
174 443
5 1 8 0 0 8320 0 7 21 0 0 6
409 121
437 121
437 503
276 503
276 441
287 441
4 2 9 0 0 4224 0 23 18 0 0 4
313 282
344 282
344 292
358 292
4 3 10 0 0 4224 0 22 18 0 0 4
313 316
345 316
345 301
358 301
4 4 11 0 0 4224 0 8 18 0 0 3
313 351
358 351
358 310
4 1 12 0 0 4224 0 25 18 0 0 3
313 246
358 246
358 283
3 0 13 0 0 4096 0 8 0 0 49 2
268 360
39 360
1 0 14 0 0 4096 0 17 0 0 48 2
204 351
68 351
2 2 15 0 0 4224 0 8 17 0 0 2
268 351
240 351
1 0 5 0 0 0 0 8 0 0 51 2
268 342
119 342
3 0 13 0 0 0 0 22 0 0 49 2
268 325
39 325
2 0 14 0 0 4096 0 22 0 0 48 2
268 316
68 316
1 0 6 0 0 0 0 22 0 0 50 2
268 307
97 307
3 0 14 0 0 0 0 23 0 0 48 2
268 291
68 291
1 0 13 0 0 0 0 6 0 0 49 2
207 282
39 282
2 2 16 0 0 4224 0 6 23 0 0 2
243 282
268 282
1 0 5 0 0 0 0 15 0 0 51 2
171 273
119 273
1 2 17 0 0 4224 0 23 15 0 0 2
268 273
207 273
1 0 14 0 0 0 0 12 0 0 48 2
206 255
68 255
3 2 18 0 0 4224 0 25 12 0 0 2
268 255
242 255
1 0 13 0 0 0 0 14 0 0 49 2
168 246
39 246
2 2 19 0 0 4224 0 25 14 0 0 2
268 246
204 246
1 0 6 0 0 0 0 25 0 0 50 2
268 237
97 237
3 2 20 0 0 4224 0 11 7 0 0 4
313 104
347 104
347 117
359 117
3 3 21 0 0 4224 0 10 7 0 0 4
313 144
348 144
348 126
359 126
4 4 22 0 0 4224 0 24 7 0 0 3
313 181
359 181
359 135
4 1 23 0 0 4224 0 9 7 0 0 3
312 65
359 65
359 108
3 0 14 0 0 0 0 24 0 0 48 2
268 190
68 190
2 0 13 0 0 0 0 24 0 0 49 2
268 181
39 181
1 0 6 0 0 0 0 24 0 0 50 2
268 172
97 172
2 0 14 0 0 0 0 10 0 0 48 2
268 153
68 153
1 0 5 0 0 0 0 10 0 0 51 2
268 135
119 135
2 2 24 0 0 4224 0 13 11 0 0 2
231 113
268 113
1 0 5 0 0 0 0 11 0 0 51 2
268 95
119 95
0 1 13 0 0 0 0 0 13 49 0 2
39 113
195 113
0 3 13 0 0 0 0 0 9 49 0 2
39 74
267 74
0 2 5 0 0 0 0 0 9 51 0 2
119 65
267 65
2 1 25 0 0 4224 0 16 9 0 0 2
230 56
267 56
0 1 6 0 0 0 0 0 16 50 0 2
97 56
194 56
1 0 14 0 0 4224 0 1 0 0 0 2
68 39
68 580
1 0 13 0 0 4224 0 2 0 0 0 2
39 39
39 579
0 0 6 0 0 4224 0 0 0 0 0 2
97 33
97 580
0 0 5 0 0 4224 0 0 0 0 0 2
119 33
119 580
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
