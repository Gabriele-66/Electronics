CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
157 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
325 176 438 273
42991634 0
0
6 Title:
5 Name:
0
0
0
26
2 +V
167 54 396 0 1 3
0 3
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
43204.9 22
0
4 LED~
171 734 235 0 2 2
10 17 18
0
0 0 112 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
391 0 0
2
43204.9 21
0
14 NO PushButton~
191 142 172 0 2 5
0 9 2
0
0 0 5232 90
0
2 S3
15 -6 29 2
6 avanti
-52 -23 -10 -15
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3124 0 0
2
43204.9 20
0
14 NO PushButton~
191 46 514 0 2 5
0 6 2
0
0 0 5232 90
0
2 S2
15 -5 29 3
4 stop
-39 -21 -11 -13
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3421 0 0
2
43204.9 19
0
14 NO PushButton~
191 84 349 0 2 5
0 10 2
0
0 0 5232 90
0
2 S1
15 -5 29 3
8 indietro
-59 -25 -3 -17
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8157 0 0
2
43204.9 18
0
7 Ground~
168 150 218 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
43204.9 17
0
7 Ground~
168 54 562 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
43204.9 16
0
7 Ground~
168 92 397 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
43204.9 15
0
2 +V
167 92 210 0 1 3
0 19
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
43204.9 14
0
2 +V
167 150 20 0 1 3
0 20
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
43204.9 13
0
2 +V
167 733 74 0 1 3
0 16
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
43204.9 12
0
2 +V
167 734 194 0 1 3
0 17
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
43204.9 11
0
5 4011~
219 286 135 0 3 22
0 9 8 7
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 2 0
1 U
3536 0 0
2
43204.9 10
0
5 4011~
219 287 252 0 3 22
0 7 6 8
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
4597 0 0
2
43204.9 9
0
5 4011~
219 287 323 0 3 22
0 10 11 12
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 3 0
1 U
3835 0 0
2
43204.9 8
0
5 4011~
219 284 403 0 3 22
0 12 6 11
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
3670 0 0
2
43204.9 7
0
5 4011~
219 416 152 0 3 22
0 7 5 4
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
5616 0 0
2
43204.9 6
0
5 4011~
219 418 266 0 3 22
0 4 12 5
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 4 0
1 U
9323 0 0
2
43204.9 5
0
5 4011~
219 556 151 0 3 22
0 4 4 14
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 4 0
1 U
317 0 0
2
43204.9 4
0
5 4011~
219 554 266 0 3 22
0 5 5 13
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 4 0
1 U
3108 0 0
2
43204.9 3
0
5 4011~
219 682 151 0 3 22
0 14 14 15
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
43204.9 2
0
5 4011~
219 687 267 0 3 22
0 13 13 18
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
43204.9 1
0
4 LED~
171 733 120 0 2 2
12 16 15
0
0 0 112 0
4 LED2
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7876 0 0
2
43204.9 0
0
9 Resistor~
219 54 450 0 4 5
0 6 3 0 1
0
0 0 112 90
3 22K
6 0 27 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
43204.9 25
0
9 Resistor~
219 150 93 0 4 5
0 9 20 0 1
0
0 0 112 90
3 22K
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
43204.9 24
0
9 Resistor~
219 92 276 0 4 5
0 10 19 0 1
0
0 0 112 90
3 22K
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
43204.9 23
0
33
2 1 3 0 0 4240 0 24 1 0 0 2
54 432
54 405
1 0 4 0 0 12432 0 18 0 0 5 5
394 257
358 257
358 194
459 194
459 152
2 0 5 0 0 12432 0 17 0 0 4 5
392 161
382 161
382 215
461 215
461 266
3 0 5 0 0 16 0 18 0 0 6 2
445 266
524 266
3 0 4 0 0 16 0 17 0 0 7 4
443 152
519 152
519 153
524 153
1 2 5 0 0 16 0 20 20 0 0 4
530 257
524 257
524 275
530 275
1 2 4 0 0 16 0 19 19 0 0 4
532 142
524 142
524 160
532 160
2 0 6 0 0 4112 0 16 0 0 9 2
260 412
199 412
2 0 6 0 0 8336 0 14 0 0 27 4
263 261
199 261
199 475
54 475
0 1 7 0 0 8336 0 0 14 11 0 5
336 135
336 179
221 179
221 243
263 243
3 1 7 0 0 16 0 13 17 0 0 4
313 135
383 135
383 143
392 143
2 3 8 0 0 12432 0 13 14 0 0 6
262 144
255 144
255 192
342 192
342 252
314 252
1 0 9 0 0 4240 0 13 0 0 32 2
262 126
150 126
1 0 10 0 0 4240 0 15 0 0 29 2
263 314
92 314
3 2 11 0 0 12432 0 16 15 0 0 6
311 403
326 403
326 357
224 357
224 332
263 332
0 1 12 0 0 8336 0 0 16 17 0 5
337 323
337 371
224 371
224 394
260 394
3 2 12 0 0 16 0 15 18 0 0 4
314 323
386 323
386 275
394 275
3 0 13 0 0 4240 0 20 0 0 19 2
581 266
657 266
1 2 13 0 0 16 0 22 22 0 0 4
663 258
657 258
657 276
663 276
3 0 14 0 0 4240 0 19 0 0 21 2
583 151
651 151
1 2 14 0 0 16 0 21 21 0 0 4
658 142
651 142
651 160
658 160
3 2 15 0 0 4240 0 21 23 0 0 3
709 151
733 151
733 130
1 1 16 0 0 4240 0 11 23 0 0 2
733 83
733 110
1 1 17 0 0 4240 0 12 2 0 0 2
734 203
734 225
3 2 18 0 0 8336 0 22 2 0 0 3
714 267
734 267
734 245
2 1 2 0 0 4240 0 4 7 0 0 2
54 531
54 556
1 1 6 0 0 16 0 24 4 0 0 2
54 468
54 497
2 1 2 0 0 16 0 5 8 0 0 2
92 366
92 391
1 1 10 0 0 16 0 26 5 0 0 2
92 294
92 332
1 2 19 0 0 4240 0 9 26 0 0 2
92 219
92 258
2 1 2 0 0 16 0 3 6 0 0 2
150 189
150 212
1 1 9 0 0 16 0 25 3 0 0 2
150 111
150 155
1 2 20 0 0 4240 0 10 25 0 0 2
150 29
150 75
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
