CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1325 608
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
17
4 LED~
171 305 225 0 1 2
10 8
0
0 0 368 90
6 GUASTO
-19 -21 23 -13
2 D3
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5130 0 0
2
43072.7 0
0
5 4049~
219 253 226 0 2 22
0 7 10
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
391 0 0
2
43072.7 0
0
5 4011~
219 199 226 0 3 22
0 10 6 11
0
0 0 96 0
4 4011
-7 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 9 0
1 U
3124 0 0
2
43072.7 0
0
4 LED~
171 303 153 0 1 2
10 8
0
0 0 368 90
9 DIREZIONE
-29 -21 34 -13
2 D2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3421 0 0
2
43072.7 0
0
5 4049~
219 152 154 0 2 22
0 7 10
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
8157 0 0
2
43072.7 0
0
5 4049~
219 151 49 0 2 22
0 7 10
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
5572 0 0
2
43072.7 11
0
5 4049~
219 138 114 0 2 22
0 3 12
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
8901 0 0
2
43072.7 10
0
7 Ground~
168 371 282 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
43072.7 9
0
4 LED~
171 302 79 0 1 2
10 8
0
0 0 368 90
6 MOTORE
-19 -21 23 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4747 0 0
2
43072.7 8
0
5 4011~
219 198 58 0 3 22
0 10 6 11
0
0 0 96 0
4 4011
-7 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 9 0
1 U
972 0 0
2
43072.7 7
0
5 4023~
219 199 105 0 4 22
0 5 4 12 9
0
0 0 96 0
4 4023
-14 -28 14 -20
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 10 0
1 U
3472 0 0
2
43072.7 6
0
5 4011~
219 263 80 0 3 22
0 11 9 8
0
0 0 96 0
4 4011
-7 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 9 0
1 U
9998 0 0
2
43072.7 5
0
5 4049~
219 154 96 0 2 22
0 6 5
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
3536 0 0
2
43072.7 4
0
13 Logic Switch~
5 123 29 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21600 270
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
1 I
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
43072.7 3
0
13 Logic Switch~
5 90 30 0 1 11
0 7
0
0 0 21728 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
1 S
-3 -26 4 -18
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
43072.7 2
0
13 Logic Switch~
5 19 30 0 1 11
0 6
0
0 0 21728 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
1 A
-3 -26 4 -18
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
43072.7 1
0
13 Logic Switch~
5 52 29 0 1 11
0 4
0
0 0 21728 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
1 C
-3 -26 4 -18
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
43072.7 0
0
24
2 0 0 0 0 0 0 1 0 0 10 2
318 226
371 226
2 0 0 0 0 0 0 4 0 0 10 2
316 154
371 154
2 1 0 0 0 0 0 2 1 0 0 2
274 226
298 226
3 1 0 0 0 0 0 3 2 0 0 2
226 226
238 226
2 0 0 0 0 0 0 3 0 0 21 2
175 235
123 235
1 0 0 0 0 0 0 3 0 0 22 2
175 217
90 217
2 1 0 0 0 0 0 5 4 0 0 2
173 154
296 154
1 0 0 0 0 0 0 5 0 0 24 2
137 154
19 154
1 3 0 0 0 0 0 9 12 0 0 2
295 80
290 80
2 1 0 0 0 0 0 9 8 0 0 3
315 80
371 80
371 276
4 2 0 0 0 0 0 11 12 0 0 4
226 105
231 105
231 89
239 89
3 1 0 0 0 0 0 10 12 0 0 4
225 58
231 58
231 71
239 71
2 3 0 0 0 0 0 7 11 0 0 2
159 114
175 114
1 0 0 0 0 0 0 7 0 0 21 2
123 114
123 113
1 2 0 0 0 0 0 11 13 0 0 2
175 96
175 96
2 1 0 0 0 0 0 6 10 0 0 2
172 49
174 49
0 2 4 0 0 0 0 0 11 23 0 2
52 105
175 105
0 1 6 0 0 0 0 0 13 24 0 2
19 96
139 96
0 2 6 0 0 0 0 0 10 24 0 2
19 67
174 67
0 1 7 0 0 0 0 0 6 22 0 2
90 49
136 49
1 0 3 0 0 0 0 14 0 0 0 2
123 41
123 426
1 0 7 0 0 0 0 15 0 0 0 2
90 42
90 425
1 0 4 0 0 0 0 17 0 0 0 2
52 41
52 426
1 0 6 0 0 0 0 16 0 0 0 2
19 42
19 426
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
