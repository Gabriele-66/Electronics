CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 90 10
176 79 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
28
10 Capacitor~
219 812 454 0 2 5
0 2 6
0
0 0 848 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3217 0 0
2
43150.7 3
0
7 Ground~
168 812 514 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3965 0 0
2
43150.7 2
0
2 +V
167 812 349 0 1 3
0 9
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8239 0 0
2
43150.7 1
0
14 NO PushButton~
191 896 456 0 2 5
0 2 6
0
0 0 4720 270
0
2 S1
14 -4 28 4
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
828 0 0
2
43150.7 0
0
10 2-In NAND~
219 218 482 0 3 22
0 15 4 10
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6187 0 0
2
5.89835e-315 0
0
10 2-In NAND~
219 246 311 0 3 22
0 14 15 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7107 0 0
2
5.89835e-315 0
0
10 2-In NAND~
219 599 429 0 3 22
0 7 8 12
0
0 0 624 692
4 7400
-7 -24 21 -16
3 U6B
-14 -27 7 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6433 0 0
2
5.89835e-315 0
0
10 2-In NAND~
219 647 384 0 3 22
0 12 6 5
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U6A
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8559 0 0
2
5.89835e-315 0
0
2 +V
167 560 585 0 1 3
0 3
0
0 0 53488 180
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
43150.7 0
0
7 Ground~
168 669 551 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5697 0 0
2
43150.7 1
0
6 74LS90
107 566 505 0 10 21
0 2 2 5 3 10 17 34 7 8
17
0
0 0 4848 602
6 74LS90
-21 -51 21 -43
2 U3
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3805 0 0
2
43150.7 2
0
9 Inverter~
13 123 384 0 2 22
0 4 14
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5219 0 0
2
43150.7 6
0
9 Inverter~
13 61 316 0 2 22
0 10 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3795 0 0
2
43150.7 7
0
4 LED~
171 593 69 0 2 2
10 4 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D8
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3637 0 0
2
43150.7 8
0
4 LED~
171 538 69 0 2 2
10 27 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D7
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3226 0 0
2
43150.7 9
0
4 LED~
171 483 73 0 2 2
10 28 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D6
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6966 0 0
2
43150.7 10
0
4 LED~
171 426 73 0 2 2
10 29 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D5
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9796 0 0
2
43150.7 11
0
4 LED~
171 368 75 0 2 2
10 33 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D4
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5952 0 0
2
43150.7 12
0
4 LED~
171 310 77 0 2 2
10 30 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D3
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3649 0 0
2
43150.7 13
0
4 LED~
171 248 77 0 2 2
10 31 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D2
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3716 0 0
2
43150.7 14
0
4 LED~
171 195 76 0 2 2
10 32 2
0
0 0 864 180
4 LED1
16 0 44 8
2 D1
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4797 0 0
2
43150.7 15
0
7 Ground~
168 657 67 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4681 0 0
2
43150.7 16
0
7 74LS244
143 389 171 0 18 37
0 19 20 21 22 23 24 25 26 4
27 28 29 33 30 31 32 13 13
0
0 0 4848 602
7 74LS244
-24 -60 25 -52
2 U1
54 -6 68 2
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
9730 0 0
2
43150.7 17
0
9 Inverter~
13 445 332 0 2 22
0 5 16
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U5A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9874 0 0
2
43150.7 18
0
2 +V
167 462 297 0 1 3
0 18
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
364 0 0
2
43150.7 20
0
7 Pulser~
4 269 413 0 10 12
0 35 36 15 37 0 0 5 5 5
8
0
0 0 4656 512
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3656 0 0
2
43150.7 21
0
7 74LS164
127 384 262 0 12 25
0 18 18 11 16 19 20 21 22 23
24 25 26
0
0 0 4848 602
7 74LS164
-24 -51 25 -43
2 U2
45 -6 59 2
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3131 0 0
2
43150.7 22
0
9 Resistor~
219 812 400 0 4 5
0 6 9 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6772 0 0
2
43150.7 4
0
52
1 4 3 0 0 4224 0 9 11 0 0 2
560 570
560 531
2 0 4 0 0 4096 0 5 0 0 3 2
194 491
126 491
0 1 4 0 0 12416 0 0 12 37 0 5
595 126
990 126
990 622
126 622
126 402
3 0 5 0 0 4096 0 8 0 0 5 2
649 357
649 332
3 1 5 0 0 16512 0 11 24 0 0 5
569 531
569 598
932 598
932 332
466 332
0 2 6 0 0 4224 0 0 8 10 0 3
812 426
658 426
658 408
1 8 7 0 0 8320 0 7 11 0 0 3
575 438
569 438
569 467
9 2 8 0 0 4224 0 11 7 0 0 3
551 467
551 420
575 420
0 1 2 0 0 4096 0 0 4 11 0 3
812 491
887 491
887 474
0 2 6 0 0 0 0 0 4 13 0 3
812 426
887 426
887 440
1 1 2 0 0 0 0 2 1 0 0 2
812 508
812 463
1 2 9 0 0 4224 0 3 28 0 0 2
812 358
812 382
1 2 6 0 0 0 0 28 1 0 0 2
812 418
812 445
3 0 10 0 0 8192 0 5 0 0 19 3
245 482
266 482
266 553
3 3 11 0 0 8320 0 27 6 0 0 3
383 293
383 311
273 311
3 1 12 0 0 8320 0 7 8 0 0 3
626 429
640 429
640 408
0 2 13 0 0 4224 0 0 13 18 0 3
380 212
64 212
64 298
17 18 13 0 0 0 0 23 23 0 0 4
424 208
424 212
379 212
379 208
5 1 10 0 0 8320 0 11 13 0 0 4
542 537
542 553
64 553
64 334
2 1 14 0 0 8320 0 12 6 0 0 3
126 366
126 302
222 302
3 0 15 0 0 4096 0 26 0 0 22 4
245 404
201 404
201 405
186 405
2 1 15 0 0 8320 0 6 5 0 0 4
222 320
186 320
186 473
194 473
4 2 16 0 0 8320 0 27 24 0 0 3
365 299
365 332
430 332
0 1 2 0 0 8320 0 0 10 25 0 3
587 543
587 545
669 545
2 1 2 0 0 0 0 11 11 0 0 4
578 531
578 543
587 543
587 531
10 6 17 0 0 12416 0 11 11 0 0 6
533 467
533 456
502 456
502 543
533 543
533 537
0 1 18 0 0 4224 0 0 25 28 0 3
410 305
462 305
462 306
2 1 18 0 0 0 0 27 27 0 0 4
401 293
401 305
410 305
410 293
1 5 19 0 0 4224 0 23 27 0 0 4
415 202
415 223
410 223
410 229
2 6 20 0 0 4224 0 23 27 0 0 4
406 202
406 222
401 222
401 229
3 7 21 0 0 4224 0 23 27 0 0 4
397 202
397 222
392 222
392 229
4 8 22 0 0 4224 0 23 27 0 0 4
388 202
388 221
383 221
383 229
5 9 23 0 0 4224 0 23 27 0 0 4
370 202
370 221
374 221
374 229
6 10 24 0 0 4224 0 23 27 0 0 4
361 202
361 221
365 221
365 229
7 11 25 0 0 4224 0 23 27 0 0 4
352 202
352 221
356 221
356 229
8 12 26 0 0 4224 0 23 27 0 0 4
343 202
343 222
347 222
347 229
1 9 4 0 0 0 0 14 23 0 0 4
595 79
595 127
415 127
415 138
1 10 27 0 0 8320 0 15 23 0 0 4
540 79
540 120
406 120
406 138
1 11 28 0 0 8320 0 16 23 0 0 4
485 83
485 112
397 112
397 138
1 12 29 0 0 8320 0 17 23 0 0 4
428 83
428 103
388 103
388 138
1 14 30 0 0 8320 0 19 23 0 0 4
312 87
312 103
361 103
361 138
1 15 31 0 0 8320 0 20 23 0 0 4
250 87
250 111
352 111
352 138
1 16 32 0 0 8320 0 21 23 0 0 4
197 86
197 119
343 119
343 138
1 13 33 0 0 4224 0 18 23 0 0 2
370 85
370 138
0 1 2 0 0 0 0 0 22 46 0 3
595 45
657 45
657 61
0 2 2 0 0 0 0 0 14 47 0 3
540 45
595 45
595 59
0 2 2 0 0 0 0 0 15 48 0 3
485 45
540 45
540 59
0 2 2 0 0 0 0 0 16 49 0 3
427 45
485 45
485 63
0 2 2 0 0 0 0 0 17 50 0 3
370 45
428 45
428 63
0 2 2 0 0 0 0 0 18 51 0 3
312 45
370 45
370 65
0 2 2 0 0 0 0 0 19 52 0 3
248 45
312 45
312 67
2 2 2 0 0 0 0 21 20 0 0 4
197 66
197 45
250 45
250 67
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
