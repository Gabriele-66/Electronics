CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 80 1313 661
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 262 331 0 1 11
0 4
0
0 0 21616 270
2 0V
11 0 25 8
2 V1
11 -10 25 -2
6 preset
-20 -22 22 -14
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4299 0 0
2
43030.7 0
0
13 Logic Switch~
5 204 321 0 1 11
0 5
0
0 0 21616 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
5 clock
-17 15 18 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
43030.7 1
0
13 Logic Switch~
5 264 193 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21616 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
8 lap test
-28 15 28 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7876 0 0
2
43030.7 2
0
13 Logic Switch~
5 351 336 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
11 0 25 8
2 V2
11 -10 25 -2
13 99 a 0/0 a 99
-47 -23 44 -15
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
43030.7 3
0
7 Ground~
168 168 288 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
43030.7 4
0
7 Ground~
168 386 288 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7100 0 0
2
43030.7 5
0
7 Ground~
168 110 286 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
43030.7 6
0
9 CC 7-Seg~
183 123 51 0 17 19
10 31 30 29 25 28 27 26 32 2
1 1 1 1 1 1 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7678 0 0
2
43030.7 7
0
7 Ground~
168 435 297 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
43030.7 8
0
7 Ground~
168 132 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
43030.7 9
0
2 +V
167 418 202 0 1 3
0 8
0
0 0 53360 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
43030.7 10
0
2 +V
167 141 202 0 1 3
0 9
0
0 0 53360 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
43030.7 11
0
7 Ground~
168 409 205 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8885 0 0
2
43030.7 12
0
9 CC 7-Seg~
183 400 53 0 17 19
10 20 19 18 14 17 16 15 33 2
1 1 1 1 1 1 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3780 0 0
2
43030.7 13
0
4 4511
219 400 157 0 14 29
0 13 12 11 10 2 8 6 15 16
17 14 18 19 20
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
9265 0 0
2
43030.7 14
0
4 4029
219 411 245 0 14 29
0 3 2 2 3 4 5 2 2 3
7 10 11 12 13
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
43030.7 15
0
7 Ground~
168 358 36 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9424 0 0
2
43030.7 16
0
7 Ground~
168 164 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9968 0 0
2
43030.7 17
0
4 4029
219 134 246 0 14 29
0 3 2 2 3 4 5 7 2 3
34 21 22 23 24
0
0 0 4336 90
4 4029
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 13 12 4 1 15 5 9 10
7 6 11 14 2 3 13 12 4 1
15 5 9 10 7 6 11 14 2 0
65 0 0 512 1 0 0 0
1 U
9281 0 0
2
5.8982e-315 0
0
4 4511
219 123 158 0 14 29
0 24 23 22 21 2 9 6 26 27
28 25 29 30 31
0
0 0 4336 90
4 4511
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8464 0 0
2
5.8982e-315 5.26354e-315
0
48
0 9 3 0 0 8192 0 0 16 17 0 3
400 372
454 372
454 279
1 0 3 0 0 0 0 4 0 0 17 2
351 348
351 372
1 0 4 0 0 4096 0 1 0 0 13 2
262 343
262 348
1 0 5 0 0 8192 0 2 0 0 5 3
205 308
205 304
225 304
6 6 5 0 0 8320 0 19 16 0 0 4
150 280
150 304
427 304
427 279
8 1 2 0 0 4096 0 19 5 0 0 4
168 280
168 284
168 284
168 282
3 1 2 0 0 0 0 19 7 0 0 2
114 280
110 280
2 1 2 0 0 4096 0 19 7 0 0 2
105 280
110 280
1 0 6 0 0 4096 0 3 0 0 10 4
265 180
267 180
267 180
265 180
7 7 6 0 0 8320 0 20 15 0 0 3
150 181
150 180
427 180
9 0 3 0 0 0 0 19 0 0 17 2
177 280
177 372
7 10 7 0 0 8320 0 19 16 0 0 5
159 286
159 360
471 360
471 209
418 209
5 5 4 0 0 8320 0 19 16 0 0 4
141 280
141 348
418 348
418 279
8 0 2 0 0 8192 0 16 0 0 24 3
445 279
445 287
436 287
3 1 2 0 0 0 0 16 6 0 0 3
391 279
391 282
386 282
2 1 2 0 0 0 0 16 6 0 0 3
382 279
382 282
386 282
4 1 3 0 0 8320 0 16 19 0 0 4
400 279
400 372
96 372
96 280
1 0 3 0 0 0 0 16 0 0 17 2
373 279
373 372
4 0 3 0 0 0 0 19 0 0 17 2
123 280
123 372
6 1 8 0 0 4224 0 15 11 0 0 4
418 180
418 188
418 188
418 187
5 1 2 0 0 4096 0 15 13 0 0 2
409 180
409 199
6 1 9 0 0 4224 0 20 12 0 0 4
141 181
141 189
141 189
141 187
5 1 2 0 0 0 0 20 10 0 0 2
132 181
132 197
7 1 2 0 0 0 0 16 9 0 0 4
436 285
436 287
435 287
435 291
9 1 2 0 0 8320 0 14 17 0 0 4
400 11
400 7
358 7
358 30
4 11 10 0 0 4224 0 15 16 0 0 2
400 174
400 215
3 12 11 0 0 4224 0 15 16 0 0 2
391 174
391 215
2 13 12 0 0 4224 0 15 16 0 0 2
382 174
382 215
1 14 13 0 0 4224 0 15 16 0 0 2
373 174
373 215
4 11 14 0 0 4224 0 14 15 0 0 3
397 89
397 110
400 110
7 8 15 0 0 4224 0 14 15 0 0 4
415 89
415 103
427 103
427 110
6 9 16 0 0 4224 0 14 15 0 0 4
409 89
409 108
418 108
418 110
5 10 17 0 0 4224 0 14 15 0 0 3
403 89
403 110
409 110
3 12 18 0 0 4224 0 14 15 0 0 2
391 89
391 110
2 13 19 0 0 4224 0 14 15 0 0 3
385 89
385 110
382 110
1 14 20 0 0 4224 0 14 15 0 0 3
379 89
379 110
373 110
9 1 2 0 0 0 0 8 18 0 0 4
123 9
123 6
164 6
164 22
4 11 21 0 0 4224 0 20 19 0 0 2
123 175
123 216
3 12 22 0 0 4224 0 20 19 0 0 2
114 175
114 216
2 13 23 0 0 4224 0 20 19 0 0 2
105 175
105 216
1 14 24 0 0 4224 0 20 19 0 0 2
96 175
96 216
4 11 25 0 0 4224 0 8 20 0 0 4
120 87
120 112
123 112
123 111
7 8 26 0 0 4224 0 8 20 0 0 4
138 87
138 102
150 102
150 111
6 9 27 0 0 4224 0 8 20 0 0 4
132 87
132 107
141 107
141 111
5 10 28 0 0 4224 0 8 20 0 0 4
126 87
126 112
132 112
132 111
3 12 29 0 0 4224 0 8 20 0 0 2
114 87
114 111
2 13 30 0 0 4224 0 8 20 0 0 4
108 87
108 112
105 112
105 111
1 14 31 0 0 4224 0 8 20 0 0 4
102 87
102 112
96 112
96 111
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
