CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 143 60 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
1 I
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43069.4 0
0
13 Logic Switch~
5 110 57 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 S
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43069.4 0
0
13 Logic Switch~
5 81 57 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 C
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43069.4 0
0
13 Logic Switch~
5 54 58 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21616 270
2 5V
-6 -17 8 -9
2 V1
-6 -26 8 -18
1 A
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43069.4 0
0
7 Ground~
168 392 144 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8157 0 0
2
43069.4 0
0
7 Ground~
168 395 179 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5572 0 0
2
43069.4 0
0
7 Ground~
168 391 85 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8901 0 0
2
43069.4 0
0
4 LED~
171 358 178 0 2 2
10 3 2
0
0 0 96 90
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7361 0 0
2
43069.4 0
0
4 LED~
171 359 145 0 2 2
10 4 2
0
0 0 96 90
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4747 0 0
2
43069.4 0
0
4 LED~
171 359 84 0 2 2
10 5 2
0
0 0 96 90
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
972 0 0
2
43069.4 0
0
9 Inverter~
13 181 177 0 2 22
0 10 9
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3472 0 0
2
43069.4 0
0
9 Inverter~
13 181 209 0 2 22
0 7 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
9998 0 0
2
43069.4 0
0
9 Inverter~
13 182 153 0 2 22
0 12 11
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
3536 0 0
2
43069.4 0
0
9 Inverter~
13 306 146 0 2 22
0 10 4
0
0 0 1136 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
9 DIREZIONE
118 0 181 8
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
4597 0 0
2
43069.4 0
0
5 4071~
219 306 180 0 3 22
0 14 13 3
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
6 MOTORE
122 -2 164 6
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
43069.4 0
0
5 4073~
219 246 191 0 4 22
0 9 6 8 13
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3670 0 0
2
43069.4 0
0
5 4081~
219 245 143 0 3 22
0 10 11 14
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
5616 0 0
2
43069.4 0
0
5 4081~
219 311 85 0 3 22
0 12 7 5
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
6 GUASTO
122 -4 164 4
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
9323 0 0
2
43069.4 0
0
23
1 2 2 0 0 8320 0 6 8 0 0 3
388 180
388 179
371 179
1 2 2 0 0 0 0 5 9 0 0 3
385 145
385 146
372 146
1 2 2 0 0 0 0 7 10 0 0 3
384 86
384 85
372 85
1 3 3 0 0 8320 0 8 15 0 0 3
351 179
351 180
339 180
1 2 4 0 0 4224 0 9 14 0 0 2
352 146
327 146
1 3 5 0 0 4224 0 10 18 0 0 2
352 85
332 85
0 2 6 0 0 4096 0 0 16 22 0 2
81 191
222 191
0 1 7 0 0 4096 0 0 12 20 0 2
143 209
166 209
2 3 8 0 0 4224 0 12 16 0 0 4
202 209
214 209
214 200
222 200
2 1 9 0 0 4224 0 11 16 0 0 4
202 177
214 177
214 182
222 182
0 1 10 0 0 4096 0 0 11 23 0 2
54 177
166 177
2 2 11 0 0 4224 0 13 17 0 0 4
203 153
213 153
213 152
221 152
0 1 12 0 0 4096 0 0 13 21 0 2
110 153
167 153
0 1 10 0 0 4096 0 0 17 23 0 2
54 134
221 134
4 2 13 0 0 4224 0 16 15 0 0 4
267 191
284 191
284 189
293 189
3 1 14 0 0 8320 0 17 15 0 0 4
266 143
284 143
284 171
293 171
0 1 10 0 0 12432 0 0 14 23 0 5
54 116
69 116
69 117
291 117
291 146
0 2 7 0 0 4096 0 0 18 20 0 2
143 94
287 94
0 1 12 0 0 4224 0 0 18 21 0 2
110 76
287 76
1 0 7 0 0 4224 0 1 0 0 0 2
143 72
143 225
1 0 12 0 0 0 0 2 0 0 0 2
110 69
110 223
1 0 6 0 0 4224 0 3 0 0 0 2
81 69
81 225
1 0 10 0 0 0 0 4 0 0 0 2
54 70
54 225
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
